-- Description:
-- Package for LUTS with ufixed format values.

-- Version history:
-- HB 2020-03-14: first design

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.fixed_pkg.all;

use work.gtl_pkg.all;

package ufixed_luts_pkg is

type eg_pt_lut_ufixed_array is array (0 to 2**(D_S_I_EG_V2.et_high-D_S_I_EG_V2.et_low+1)-1) of ufixed(7 downto -20);
constant EG_PT_LUT_UFIXED : eg_pt_lut_ufixed_array := (
"0000000001001100110011001100", "0000000011001100110011001100", "0000000101001100110011001100", "0000000111001100110011001100", 
"0000001001001100110011001100", "0000001011001100110011001100", "0000001101001100110011001100", "0000001111001100110011001100", 
"0000010001001100110011001100", "0000010011001100110011001100", "0000010101001100110011001100", "0000010111001100110011001100", 
"0000011001001100110011001100", "0000011011001100110011001100", "0000011101001100110011001100", "0000011111001100110011001100", 
"0000100001001100110011001100", "0000100011001100110011001100", "0000100101001100110011001100", "0000100111001100110011001100", 
"0000101001001100110011001100", "0000101011001100110011001100", "0000101101001100110011001100", "0000101111001100110011001100", 
"0000110001001100110011001100", "0000110011001100110011001100", "0000110101001100110011001100", "0000110111001100110011001100", 
"0000111001001100110011001100", "0000111011001100110011001100", "0000111101001100110011001100", "0000111111001100110011001100", 
"0001000001001100110011001100", "0001000011001100110011001100", "0001000101001100110011001100", "0001000111001100110011001100", 
"0001001001001100110011001100", "0001001011001100110011001100", "0001001101001100110011001100", "0001001111001100110011001100", 
"0001010001001100110011001100", "0001010011001100110011001100", "0001010101001100110011001100", "0001010111001100110011001100", 
"0001011001001100110011001100", "0001011011001100110011001100", "0001011101001100110011001100", "0001011111001100110011001100", 
"0001100001001100110011001100", "0001100011001100110011001100", "0001100101001100110011001100", "0001100111001100110011001100", 
"0001101001001100110011001100", "0001101011001100110011001100", "0001101101001100110011001100", "0001101111001100110011001100", 
"0001110001001100110011001100", "0001110011001100110011001100", "0001110101001100110011001100", "0001110111001100110011001100", 
"0001111001001100110011001100", "0001111011001100110011001100", "0001111101001100110011001100", "0001111111001100110011001100", 
"0010000001001100110011001100", "0010000011001100110011001100", "0010000101001100110011001100", "0010000111001100110011001100", 
"0010001001001100110011001100", "0010001011001100110011001100", "0010001101001100110011001100", "0010001111001100110011001100", 
"0010010001001100110011001100", "0010010011001100110011001100", "0010010101001100110011001100", "0010010111001100110011001100", 
"0010011001001100110011001100", "0010011011001100110011001100", "0010011101001100110011001100", "0010011111001100110011001100", 
"0010100001001100110011001100", "0010100011001100110011001100", "0010100101001100110011001100", "0010100111001100110011001100", 
"0010101001001100110011001100", "0010101011001100110011001100", "0010101101001100110011001100", "0010101111001100110011001100", 
"0010110001001100110011001100", "0010110011001100110011001100", "0010110101001100110011001100", "0010110111001100110011001100", 
"0010111001001100110011001100", "0010111011001100110011001100", "0010111101001100110011001100", "0010111111001100110011001100", 
"0011000001001100110011001100", "0011000011001100110011001100", "0011000101001100110011001100", "0011000111001100110011001100", 
"0011001001001100110011001100", "0011001011001100110011001100", "0011001101001100110011001100", "0011001111001100110011001100", 
"0011010001001100110011001100", "0011010011001100110011001100", "0011010101001100110011001100", "0011010111001100110011001100", 
"0011011001001100110011001100", "0011011011001100110011001100", "0011011101001100110011001100", "0011011111001100110011001100", 
"0011100001001100110011001100", "0011100011001100110011001100", "0011100101001100110011001100", "0011100111001100110011001100", 
"0011101001001100110011001100", "0011101011001100110011001100", "0011101101001100110011001100", "0011101111001100110011001100", 
"0011110001001100110011001100", "0011110011001100110011001100", "0011110101001100110011001100", "0011110111001100110011001100", 
"0011111001001100110011001100", "0011111011001100110011001100", "0011111101001100110011001100", "0011111111001100110011001100", 
"0100000001001100110011001100", "0100000011001100110011001100", "0100000101001100110011001100", "0100000111001100110011001100", 
"0100001001001100110011001100", "0100001011001100110011001100", "0100001101001100110011001100", "0100001111001100110011001100", 
"0100010001001100110011001100", "0100010011001100110011001100", "0100010101001100110011001100", "0100010111001100110011001100", 
"0100011001001100110011001100", "0100011011001100110011001100", "0100011101001100110011001100", "0100011111001100110011001100", 
"0100100001001100110011001100", "0100100011001100110011001100", "0100100101001100110011001100", "0100100111001100110011001100", 
"0100101001001100110011001100", "0100101011001100110011001100", "0100101101001100110011001100", "0100101111001100110011001100", 
"0100110001001100110011001100", "0100110011001100110011001100", "0100110101001100110011001100", "0100110111001100110011001100", 
"0100111001001100110011001100", "0100111011001100110011001100", "0100111101001100110011001100", "0100111111001100110011001100", 
"0101000001001100110011001100", "0101000011001100110011001100", "0101000101001100110011001100", "0101000111001100110011001100", 
"0101001001001100110011001100", "0101001011001100110011001100", "0101001101001100110011001100", "0101001111001100110011001100", 
"0101010001001100110011001100", "0101010011001100110011001100", "0101010101001100110011001100", "0101010111001100110011001100", 
"0101011001001100110011001100", "0101011011001100110011001100", "0101011101001100110011001100", "0101011111001100110011001100", 
"0101100001001100110011001100", "0101100011001100110011001100", "0101100101001100110011001100", "0101100111001100110011001100", 
"0101101001001100110011001100", "0101101011001100110011001100", "0101101101001100110011001100", "0101101111001100110011001100", 
"0101110001001100110011001100", "0101110011001100110011001100", "0101110101001100110011001100", "0101110111001100110011001100", 
"0101111001001100110011001100", "0101111011001100110011001100", "0101111101001100110011001100", "0101111111001100110011001100", 
"0110000001001100110011001100", "0110000011001100110011001100", "0110000101001100110011001100", "0110000111001100110011001100", 
"0110001001001100110011001100", "0110001011001100110011001100", "0110001101001100110011001100", "0110001111001100110011001100", 
"0110010001001100110011001100", "0110010011001100110011001100", "0110010101001100110011001100", "0110010111001100110011001100", 
"0110011001001100110011001100", "0110011011001100110011001100", "0110011101001100110011001100", "0110011111001100110011001100", 
"0110100001001100110011001100", "0110100011001100110011001100", "0110100101001100110011001100", "0110100111001100110011001100", 
"0110101001001100110011001100", "0110101011001100110011001100", "0110101101001100110011001100", "0110101111001100110011001100", 
"0110110001001100110011001100", "0110110011001100110011001100", "0110110101001100110011001100", "0110110111001100110011001100", 
"0110111001001100110011001100", "0110111011001100110011001100", "0110111101001100110011001100", "0110111111001100110011001100", 
"0111000001001100110011001100", "0111000011001100110011001100", "0111000101001100110011001100", "0111000111001100110011001100", 
"0111001001001100110011001100", "0111001011001100110011001100", "0111001101001100110011001100", "0111001111001100110011001100", 
"0111010001001100110011001100", "0111010011001100110011001100", "0111010101001100110011001100", "0111010111001100110011001100", 
"0111011001001100110011001100", "0111011011001100110011001100", "0111011101001100110011001100", "0111011111001100110011001100", 
"0111100001001100110011001100", "0111100011001100110011001100", "0111100101001100110011001100", "0111100111001100110011001100", 
"0111101001001100110011001100", "0111101011001100110011001100", "0111101101001100110011001100", "0111101111001100110011001100", 
"0111110001001100110011001100", "0111110011001100110011001100", "0111110101001100110011001100", "0111110111001100110011001100", 
"0111111001001100110011001100", "0111111011001100110011001100", "0111111101001100110011001100", "0111111111001100110011001100", 
"1000000001001100110011001100", "1000000011001100110011001100", "1000000101001100110011001100", "1000000111001100110011001100", 
"1000001001001100110011001100", "1000001011001100110011001100", "1000001101001100110011001100", "1000001111001100110011001100", 
"1000010001001100110011001100", "1000010011001100110011001100", "1000010101001100110011001100", "1000010111001100110011001100", 
"1000011001001100110011001100", "1000011011001100110011001100", "1000011101001100110011001100", "1000011111001100110011001100", 
"1000100001001100110011001100", "1000100011001100110011001100", "1000100101001100110011001100", "1000100111001100110011001100", 
"1000101001001100110011001100", "1000101011001100110011001100", "1000101101001100110011001100", "1000101111001100110011001100", 
"1000110001001100110011001100", "1000110011001100110011001100", "1000110101001100110011001100", "1000110111001100110011001100", 
"1000111001001100110011001100", "1000111011001100110011001100", "1000111101001100110011001100", "1000111111001100110011001100", 
"1001000001001100110011001100", "1001000011001100110011001100", "1001000101001100110011001100", "1001000111001100110011001100", 
"1001001001001100110011001100", "1001001011001100110011001100", "1001001101001100110011001100", "1001001111001100110011001100", 
"1001010001001100110011001100", "1001010011001100110011001100", "1001010101001100110011001100", "1001010111001100110011001100", 
"1001011001001100110011001100", "1001011011001100110011001100", "1001011101001100110011001100", "1001011111001100110011001100", 
"1001100001001100110011001100", "1001100011001100110011001100", "1001100101001100110011001100", "1001100111001100110011001100", 
"1001101001001100110011001100", "1001101011001100110011001100", "1001101101001100110011001100", "1001101111001100110011001100", 
"1001110001001100110011001100", "1001110011001100110011001100", "1001110101001100110011001100", "1001110111001100110011001100", 
"1001111001001100110011001100", "1001111011001100110011001100", "1001111101001100110011001100", "1001111111001100110011001100", 
"1010000001001100110011001100", "1010000011001100110011001100", "1010000101001100110011001100", "1010000111001100110011001100", 
"1010001001001100110011001100", "1010001011001100110011001100", "1010001101001100110011001100", "1010001111001100110011001100", 
"1010010001001100110011001100", "1010010011001100110011001100", "1010010101001100110011001100", "1010010111001100110011001100", 
"1010011001001100110011001100", "1010011011001100110011001100", "1010011101001100110011001100", "1010011111001100110011001100", 
"1010100001001100110011001100", "1010100011001100110011001100", "1010100101001100110011001100", "1010100111001100110011001100", 
"1010101001001100110011001100", "1010101011001100110011001100", "1010101101001100110011001100", "1010101111001100110011001100", 
"1010110001001100110011001100", "1010110011001100110011001100", "1010110101001100110011001100", "1010110111001100110011001100", 
"1010111001001100110011001100", "1010111011001100110011001100", "1010111101001100110011001100", "1010111111001100110011001100", 
"1011000001001100110011001100", "1011000011001100110011001100", "1011000101001100110011001100", "1011000111001100110011001100", 
"1011001001001100110011001100", "1011001011001100110011001100", "1011001101001100110011001100", "1011001111001100110011001100", 
"1011010001001100110011001100", "1011010011001100110011001100", "1011010101001100110011001100", "1011010111001100110011001100", 
"1011011001001100110011001100", "1011011011001100110011001100", "1011011101001100110011001100", "1011011111001100110011001100", 
"1011100001001100110011001100", "1011100011001100110011001100", "1011100101001100110011001100", "1011100111001100110011001100", 
"1011101001001100110011001100", "1011101011001100110011001100", "1011101101001100110011001100", "1011101111001100110011001100", 
"1011110001001100110011001100", "1011110011001100110011001100", "1011110101001100110011001100", "1011110111001100110011001100", 
"1011111001001100110011001100", "1011111011001100110011001100", "1011111101001100110011001100", "1011111111001100110011001100", 
"1100000001001100110011001100", "1100000011001100110011001100", "1100000101001100110011001100", "1100000111001100110011001100", 
"1100001001001100110011001100", "1100001011001100110011001100", "1100001101001100110011001100", "1100001111001100110011001100", 
"1100010001001100110011001100", "1100010011001100110011001100", "1100010101001100110011001100", "1100010111001100110011001100", 
"1100011001001100110011001100", "1100011011001100110011001100", "1100011101001100110011001100", "1100011111001100110011001100", 
"1100100001001100110011001100", "1100100011001100110011001100", "1100100101001100110011001100", "1100100111001100110011001100", 
"1100101001001100110011001100", "1100101011001100110011001100", "1100101101001100110011001100", "1100101111001100110011001100", 
"1100110001001100110011001100", "1100110011001100110011001100", "1100110101001100110011001100", "1100110111001100110011001100", 
"1100111001001100110011001100", "1100111011001100110011001100", "1100111101001100110011001100", "1100111111001100110011001100", 
"1101000001001100110011001100", "1101000011001100110011001100", "1101000101001100110011001100", "1101000111001100110011001100", 
"1101001001001100110011001100", "1101001011001100110011001100", "1101001101001100110011001100", "1101001111001100110011001100", 
"1101010001001100110011001100", "1101010011001100110011001100", "1101010101001100110011001100", "1101010111001100110011001100", 
"1101011001001100110011001100", "1101011011001100110011001100", "1101011101001100110011001100", "1101011111001100110011001100", 
"1101100001001100110011001100", "1101100011001100110011001100", "1101100101001100110011001100", "1101100111001100110011001100", 
"1101101001001100110011001100", "1101101011001100110011001100", "1101101101001100110011001100", "1101101111001100110011001100", 
"1101110001001100110011001100", "1101110011001100110011001100", "1101110101001100110011001100", "1101110111001100110011001100", 
"1101111001001100110011001100", "1101111011001100110011001100", "1101111101001100110011001100", "1101111111001100110011001100", 
"1110000001001100110011001100", "1110000011001100110011001100", "1110000101001100110011001100", "1110000111001100110011001100", 
"1110001001001100110011001100", "1110001011001100110011001100", "1110001101001100110011001100", "1110001111001100110011001100", 
"1110010001001100110011001100", "1110010011001100110011001100", "1110010101001100110011001100", "1110010111001100110011001100", 
"1110011001001100110011001100", "1110011011001100110011001100", "1110011101001100110011001100", "1110011111001100110011001100", 
"1110100001001100110011001100", "1110100011001100110011001100", "1110100101001100110011001100", "1110100111001100110011001100", 
"1110101001001100110011001100", "1110101011001100110011001100", "1110101101001100110011001100", "1110101111001100110011001100", 
"1110110001001100110011001100", "1110110011001100110011001100", "1110110101001100110011001100", "1110110111001100110011001100", 
"1110111001001100110011001100", "1110111011001100110011001100", "1110111101001100110011001100", "1110111111001100110011001100", 
"1111000001001100110011001100", "1111000011001100110011001100", "1111000101001100110011001100", "1111000111001100110011001100", 
"1111001001001100110011001100", "1111001011001100110011001100", "1111001101001100110011001100", "1111001111001100110011001100", 
"1111010001001100110011001100", "1111010011001100110011001100", "1111010101001100110011001100", "1111010111001100110011001100", 
"1111011001001100110011001100", "1111011011001100110011001100", "1111011101001100110011001100", "1111011111001100110011001100", 
"1111100001001100110011001100", "1111100011001100110011001100", "1111100101001100110011001100", "1111100111001100110011001100", 
"1111101001001100110011001100", "1111101011001100110011001100", "1111101101001100110011001100", "1111101111001100110011001100", 
"1111110001001100110011001100", "1111110011001100110011001100", "1111110101001100110011001100", "1111110111001100110011001100", 
"1111111001001100110011001100", "1111111011001100110011001100", "1111111101001100110011001100", "1111111111001100110011001100"
);
type jet_pt_lut_ufixed_array is array (0 to 2**(D_S_I_JET_V2.et_high-D_S_I_JET_V2.et_low+1)-1) of ufixed(9 downto -20);
constant JET_PT_LUT_UFIXED : jet_pt_lut_ufixed_array := (
"000000000001001100110011001100", "000000000011001100110011001100", "000000000101001100110011001100", "000000000111001100110011001100", 
"000000001001001100110011001100", "000000001011001100110011001100", "000000001101001100110011001100", "000000001111001100110011001100", 
"000000010001001100110011001100", "000000010011001100110011001100", "000000010101001100110011001100", "000000010111001100110011001100", 
"000000011001001100110011001100", "000000011011001100110011001100", "000000011101001100110011001100", "000000011111001100110011001100", 
"000000100001001100110011001100", "000000100011001100110011001100", "000000100101001100110011001100", "000000100111001100110011001100", 
"000000101001001100110011001100", "000000101011001100110011001100", "000000101101001100110011001100", "000000101111001100110011001100", 
"000000110001001100110011001100", "000000110011001100110011001100", "000000110101001100110011001100", "000000110111001100110011001100", 
"000000111001001100110011001100", "000000111011001100110011001100", "000000111101001100110011001100", "000000111111001100110011001100", 
"000001000001001100110011001100", "000001000011001100110011001100", "000001000101001100110011001100", "000001000111001100110011001100", 
"000001001001001100110011001100", "000001001011001100110011001100", "000001001101001100110011001100", "000001001111001100110011001100", 
"000001010001001100110011001100", "000001010011001100110011001100", "000001010101001100110011001100", "000001010111001100110011001100", 
"000001011001001100110011001100", "000001011011001100110011001100", "000001011101001100110011001100", "000001011111001100110011001100", 
"000001100001001100110011001100", "000001100011001100110011001100", "000001100101001100110011001100", "000001100111001100110011001100", 
"000001101001001100110011001100", "000001101011001100110011001100", "000001101101001100110011001100", "000001101111001100110011001100", 
"000001110001001100110011001100", "000001110011001100110011001100", "000001110101001100110011001100", "000001110111001100110011001100", 
"000001111001001100110011001100", "000001111011001100110011001100", "000001111101001100110011001100", "000001111111001100110011001100", 
"000010000001001100110011001100", "000010000011001100110011001100", "000010000101001100110011001100", "000010000111001100110011001100", 
"000010001001001100110011001100", "000010001011001100110011001100", "000010001101001100110011001100", "000010001111001100110011001100", 
"000010010001001100110011001100", "000010010011001100110011001100", "000010010101001100110011001100", "000010010111001100110011001100", 
"000010011001001100110011001100", "000010011011001100110011001100", "000010011101001100110011001100", "000010011111001100110011001100", 
"000010100001001100110011001100", "000010100011001100110011001100", "000010100101001100110011001100", "000010100111001100110011001100", 
"000010101001001100110011001100", "000010101011001100110011001100", "000010101101001100110011001100", "000010101111001100110011001100", 
"000010110001001100110011001100", "000010110011001100110011001100", "000010110101001100110011001100", "000010110111001100110011001100", 
"000010111001001100110011001100", "000010111011001100110011001100", "000010111101001100110011001100", "000010111111001100110011001100", 
"000011000001001100110011001100", "000011000011001100110011001100", "000011000101001100110011001100", "000011000111001100110011001100", 
"000011001001001100110011001100", "000011001011001100110011001100", "000011001101001100110011001100", "000011001111001100110011001100", 
"000011010001001100110011001100", "000011010011001100110011001100", "000011010101001100110011001100", "000011010111001100110011001100", 
"000011011001001100110011001100", "000011011011001100110011001100", "000011011101001100110011001100", "000011011111001100110011001100", 
"000011100001001100110011001100", "000011100011001100110011001100", "000011100101001100110011001100", "000011100111001100110011001100", 
"000011101001001100110011001100", "000011101011001100110011001100", "000011101101001100110011001100", "000011101111001100110011001100", 
"000011110001001100110011001100", "000011110011001100110011001100", "000011110101001100110011001100", "000011110111001100110011001100", 
"000011111001001100110011001100", "000011111011001100110011001100", "000011111101001100110011001100", "000011111111001100110011001100", 
"000100000001001100110011001100", "000100000011001100110011001100", "000100000101001100110011001100", "000100000111001100110011001100", 
"000100001001001100110011001100", "000100001011001100110011001100", "000100001101001100110011001100", "000100001111001100110011001100", 
"000100010001001100110011001100", "000100010011001100110011001100", "000100010101001100110011001100", "000100010111001100110011001100", 
"000100011001001100110011001100", "000100011011001100110011001100", "000100011101001100110011001100", "000100011111001100110011001100", 
"000100100001001100110011001100", "000100100011001100110011001100", "000100100101001100110011001100", "000100100111001100110011001100", 
"000100101001001100110011001100", "000100101011001100110011001100", "000100101101001100110011001100", "000100101111001100110011001100", 
"000100110001001100110011001100", "000100110011001100110011001100", "000100110101001100110011001100", "000100110111001100110011001100", 
"000100111001001100110011001100", "000100111011001100110011001100", "000100111101001100110011001100", "000100111111001100110011001100", 
"000101000001001100110011001100", "000101000011001100110011001100", "000101000101001100110011001100", "000101000111001100110011001100", 
"000101001001001100110011001100", "000101001011001100110011001100", "000101001101001100110011001100", "000101001111001100110011001100", 
"000101010001001100110011001100", "000101010011001100110011001100", "000101010101001100110011001100", "000101010111001100110011001100", 
"000101011001001100110011001100", "000101011011001100110011001100", "000101011101001100110011001100", "000101011111001100110011001100", 
"000101100001001100110011001100", "000101100011001100110011001100", "000101100101001100110011001100", "000101100111001100110011001100", 
"000101101001001100110011001100", "000101101011001100110011001100", "000101101101001100110011001100", "000101101111001100110011001100", 
"000101110001001100110011001100", "000101110011001100110011001100", "000101110101001100110011001100", "000101110111001100110011001100", 
"000101111001001100110011001100", "000101111011001100110011001100", "000101111101001100110011001100", "000101111111001100110011001100", 
"000110000001001100110011001100", "000110000011001100110011001100", "000110000101001100110011001100", "000110000111001100110011001100", 
"000110001001001100110011001100", "000110001011001100110011001100", "000110001101001100110011001100", "000110001111001100110011001100", 
"000110010001001100110011001100", "000110010011001100110011001100", "000110010101001100110011001100", "000110010111001100110011001100", 
"000110011001001100110011001100", "000110011011001100110011001100", "000110011101001100110011001100", "000110011111001100110011001100", 
"000110100001001100110011001100", "000110100011001100110011001100", "000110100101001100110011001100", "000110100111001100110011001100", 
"000110101001001100110011001100", "000110101011001100110011001100", "000110101101001100110011001100", "000110101111001100110011001100", 
"000110110001001100110011001100", "000110110011001100110011001100", "000110110101001100110011001100", "000110110111001100110011001100", 
"000110111001001100110011001100", "000110111011001100110011001100", "000110111101001100110011001100", "000110111111001100110011001100", 
"000111000001001100110011001100", "000111000011001100110011001100", "000111000101001100110011001100", "000111000111001100110011001100", 
"000111001001001100110011001100", "000111001011001100110011001100", "000111001101001100110011001100", "000111001111001100110011001100", 
"000111010001001100110011001100", "000111010011001100110011001100", "000111010101001100110011001100", "000111010111001100110011001100", 
"000111011001001100110011001100", "000111011011001100110011001100", "000111011101001100110011001100", "000111011111001100110011001100", 
"000111100001001100110011001100", "000111100011001100110011001100", "000111100101001100110011001100", "000111100111001100110011001100", 
"000111101001001100110011001100", "000111101011001100110011001100", "000111101101001100110011001100", "000111101111001100110011001100", 
"000111110001001100110011001100", "000111110011001100110011001100", "000111110101001100110011001100", "000111110111001100110011001100", 
"000111111001001100110011001100", "000111111011001100110011001100", "000111111101001100110011001100", "000111111111001100110011001100", 
"001000000001001100110011001100", "001000000011001100110011001100", "001000000101001100110011001100", "001000000111001100110011001100", 
"001000001001001100110011001100", "001000001011001100110011001100", "001000001101001100110011001100", "001000001111001100110011001100", 
"001000010001001100110011001100", "001000010011001100110011001100", "001000010101001100110011001100", "001000010111001100110011001100", 
"001000011001001100110011001100", "001000011011001100110011001100", "001000011101001100110011001100", "001000011111001100110011001100", 
"001000100001001100110011001100", "001000100011001100110011001100", "001000100101001100110011001100", "001000100111001100110011001100", 
"001000101001001100110011001100", "001000101011001100110011001100", "001000101101001100110011001100", "001000101111001100110011001100", 
"001000110001001100110011001100", "001000110011001100110011001100", "001000110101001100110011001100", "001000110111001100110011001100", 
"001000111001001100110011001100", "001000111011001100110011001100", "001000111101001100110011001100", "001000111111001100110011001100", 
"001001000001001100110011001100", "001001000011001100110011001100", "001001000101001100110011001100", "001001000111001100110011001100", 
"001001001001001100110011001100", "001001001011001100110011001100", "001001001101001100110011001100", "001001001111001100110011001100", 
"001001010001001100110011001100", "001001010011001100110011001100", "001001010101001100110011001100", "001001010111001100110011001100", 
"001001011001001100110011001100", "001001011011001100110011001100", "001001011101001100110011001100", "001001011111001100110011001100", 
"001001100001001100110011001100", "001001100011001100110011001100", "001001100101001100110011001100", "001001100111001100110011001100", 
"001001101001001100110011001100", "001001101011001100110011001100", "001001101101001100110011001100", "001001101111001100110011001100", 
"001001110001001100110011001100", "001001110011001100110011001100", "001001110101001100110011001100", "001001110111001100110011001100", 
"001001111001001100110011001100", "001001111011001100110011001100", "001001111101001100110011001100", "001001111111001100110011001100", 
"001010000001001100110011001100", "001010000011001100110011001100", "001010000101001100110011001100", "001010000111001100110011001100", 
"001010001001001100110011001100", "001010001011001100110011001100", "001010001101001100110011001100", "001010001111001100110011001100", 
"001010010001001100110011001100", "001010010011001100110011001100", "001010010101001100110011001100", "001010010111001100110011001100", 
"001010011001001100110011001100", "001010011011001100110011001100", "001010011101001100110011001100", "001010011111001100110011001100", 
"001010100001001100110011001100", "001010100011001100110011001100", "001010100101001100110011001100", "001010100111001100110011001100", 
"001010101001001100110011001100", "001010101011001100110011001100", "001010101101001100110011001100", "001010101111001100110011001100", 
"001010110001001100110011001100", "001010110011001100110011001100", "001010110101001100110011001100", "001010110111001100110011001100", 
"001010111001001100110011001100", "001010111011001100110011001100", "001010111101001100110011001100", "001010111111001100110011001100", 
"001011000001001100110011001100", "001011000011001100110011001100", "001011000101001100110011001100", "001011000111001100110011001100", 
"001011001001001100110011001100", "001011001011001100110011001100", "001011001101001100110011001100", "001011001111001100110011001100", 
"001011010001001100110011001100", "001011010011001100110011001100", "001011010101001100110011001100", "001011010111001100110011001100", 
"001011011001001100110011001100", "001011011011001100110011001100", "001011011101001100110011001100", "001011011111001100110011001100", 
"001011100001001100110011001100", "001011100011001100110011001100", "001011100101001100110011001100", "001011100111001100110011001100", 
"001011101001001100110011001100", "001011101011001100110011001100", "001011101101001100110011001100", "001011101111001100110011001100", 
"001011110001001100110011001100", "001011110011001100110011001100", "001011110101001100110011001100", "001011110111001100110011001100", 
"001011111001001100110011001100", "001011111011001100110011001100", "001011111101001100110011001100", "001011111111001100110011001100", 
"001100000001001100110011001100", "001100000011001100110011001100", "001100000101001100110011001100", "001100000111001100110011001100", 
"001100001001001100110011001100", "001100001011001100110011001100", "001100001101001100110011001100", "001100001111001100110011001100", 
"001100010001001100110011001100", "001100010011001100110011001100", "001100010101001100110011001100", "001100010111001100110011001100", 
"001100011001001100110011001100", "001100011011001100110011001100", "001100011101001100110011001100", "001100011111001100110011001100", 
"001100100001001100110011001100", "001100100011001100110011001100", "001100100101001100110011001100", "001100100111001100110011001100", 
"001100101001001100110011001100", "001100101011001100110011001100", "001100101101001100110011001100", "001100101111001100110011001100", 
"001100110001001100110011001100", "001100110011001100110011001100", "001100110101001100110011001100", "001100110111001100110011001100", 
"001100111001001100110011001100", "001100111011001100110011001100", "001100111101001100110011001100", "001100111111001100110011001100", 
"001101000001001100110011001100", "001101000011001100110011001100", "001101000101001100110011001100", "001101000111001100110011001100", 
"001101001001001100110011001100", "001101001011001100110011001100", "001101001101001100110011001100", "001101001111001100110011001100", 
"001101010001001100110011001100", "001101010011001100110011001100", "001101010101001100110011001100", "001101010111001100110011001100", 
"001101011001001100110011001100", "001101011011001100110011001100", "001101011101001100110011001100", "001101011111001100110011001100", 
"001101100001001100110011001100", "001101100011001100110011001100", "001101100101001100110011001100", "001101100111001100110011001100", 
"001101101001001100110011001100", "001101101011001100110011001100", "001101101101001100110011001100", "001101101111001100110011001100", 
"001101110001001100110011001100", "001101110011001100110011001100", "001101110101001100110011001100", "001101110111001100110011001100", 
"001101111001001100110011001100", "001101111011001100110011001100", "001101111101001100110011001100", "001101111111001100110011001100", 
"001110000001001100110011001100", "001110000011001100110011001100", "001110000101001100110011001100", "001110000111001100110011001100", 
"001110001001001100110011001100", "001110001011001100110011001100", "001110001101001100110011001100", "001110001111001100110011001100", 
"001110010001001100110011001100", "001110010011001100110011001100", "001110010101001100110011001100", "001110010111001100110011001100", 
"001110011001001100110011001100", "001110011011001100110011001100", "001110011101001100110011001100", "001110011111001100110011001100", 
"001110100001001100110011001100", "001110100011001100110011001100", "001110100101001100110011001100", "001110100111001100110011001100", 
"001110101001001100110011001100", "001110101011001100110011001100", "001110101101001100110011001100", "001110101111001100110011001100", 
"001110110001001100110011001100", "001110110011001100110011001100", "001110110101001100110011001100", "001110110111001100110011001100", 
"001110111001001100110011001100", "001110111011001100110011001100", "001110111101001100110011001100", "001110111111001100110011001100", 
"001111000001001100110011001100", "001111000011001100110011001100", "001111000101001100110011001100", "001111000111001100110011001100", 
"001111001001001100110011001100", "001111001011001100110011001100", "001111001101001100110011001100", "001111001111001100110011001100", 
"001111010001001100110011001100", "001111010011001100110011001100", "001111010101001100110011001100", "001111010111001100110011001100", 
"001111011001001100110011001100", "001111011011001100110011001100", "001111011101001100110011001100", "001111011111001100110011001100", 
"001111100001001100110011001100", "001111100011001100110011001100", "001111100101001100110011001100", "001111100111001100110011001100", 
"001111101001001100110011001100", "001111101011001100110011001100", "001111101101001100110011001100", "001111101111001100110011001100", 
"001111110001001100110011001100", "001111110011001100110011001100", "001111110101001100110011001100", "001111110111001100110011001100", 
"001111111001001100110011001100", "001111111011001100110011001100", "001111111101001100110011001100", "001111111111001100110011001100", 
"010000000001001100110011001100", "010000000011001100110011001100", "010000000101001100110011001100", "010000000111001100110011001100", 
"010000001001001100110011001100", "010000001011001100110011001100", "010000001101001100110011001100", "010000001111001100110011001100", 
"010000010001001100110011001100", "010000010011001100110011001100", "010000010101001100110011001100", "010000010111001100110011001100", 
"010000011001001100110011001100", "010000011011001100110011001100", "010000011101001100110011001100", "010000011111001100110011001100", 
"010000100001001100110011001100", "010000100011001100110011001100", "010000100101001100110011001100", "010000100111001100110011001100", 
"010000101001001100110011001100", "010000101011001100110011001100", "010000101101001100110011001100", "010000101111001100110011001100", 
"010000110001001100110011001100", "010000110011001100110011001100", "010000110101001100110011001100", "010000110111001100110011001100", 
"010000111001001100110011001100", "010000111011001100110011001100", "010000111101001100110011001100", "010000111111001100110011001100", 
"010001000001001100110011001100", "010001000011001100110011001100", "010001000101001100110011001100", "010001000111001100110011001100", 
"010001001001001100110011001100", "010001001011001100110011001100", "010001001101001100110011001100", "010001001111001100110011001100", 
"010001010001001100110011001100", "010001010011001100110011001100", "010001010101001100110011001100", "010001010111001100110011001100", 
"010001011001001100110011001100", "010001011011001100110011001100", "010001011101001100110011001100", "010001011111001100110011001100", 
"010001100001001100110011001100", "010001100011001100110011001100", "010001100101001100110011001100", "010001100111001100110011001100", 
"010001101001001100110011001100", "010001101011001100110011001100", "010001101101001100110011001100", "010001101111001100110011001100", 
"010001110001001100110011001100", "010001110011001100110011001100", "010001110101001100110011001100", "010001110111001100110011001100", 
"010001111001001100110011001100", "010001111011001100110011001100", "010001111101001100110011001100", "010001111111001100110011001100", 
"010010000001001100110011001100", "010010000011001100110011001100", "010010000101001100110011001100", "010010000111001100110011001100", 
"010010001001001100110011001100", "010010001011001100110011001100", "010010001101001100110011001100", "010010001111001100110011001100", 
"010010010001001100110011001100", "010010010011001100110011001100", "010010010101001100110011001100", "010010010111001100110011001100", 
"010010011001001100110011001100", "010010011011001100110011001100", "010010011101001100110011001100", "010010011111001100110011001100", 
"010010100001001100110011001100", "010010100011001100110011001100", "010010100101001100110011001100", "010010100111001100110011001100", 
"010010101001001100110011001100", "010010101011001100110011001100", "010010101101001100110011001100", "010010101111001100110011001100", 
"010010110001001100110011001100", "010010110011001100110011001100", "010010110101001100110011001100", "010010110111001100110011001100", 
"010010111001001100110011001100", "010010111011001100110011001100", "010010111101001100110011001100", "010010111111001100110011001100", 
"010011000001001100110011001100", "010011000011001100110011001100", "010011000101001100110011001100", "010011000111001100110011001100", 
"010011001001001100110011001100", "010011001011001100110011001100", "010011001101001100110011001100", "010011001111001100110011001100", 
"010011010001001100110011001100", "010011010011001100110011001100", "010011010101001100110011001100", "010011010111001100110011001100", 
"010011011001001100110011001100", "010011011011001100110011001100", "010011011101001100110011001100", "010011011111001100110011001100", 
"010011100001001100110011001100", "010011100011001100110011001100", "010011100101001100110011001100", "010011100111001100110011001100", 
"010011101001001100110011001100", "010011101011001100110011001100", "010011101101001100110011001100", "010011101111001100110011001100", 
"010011110001001100110011001100", "010011110011001100110011001100", "010011110101001100110011001100", "010011110111001100110011001100", 
"010011111001001100110011001100", "010011111011001100110011001100", "010011111101001100110011001100", "010011111111001100110011001100", 
"010100000001001100110011001100", "010100000011001100110011001100", "010100000101001100110011001100", "010100000111001100110011001100", 
"010100001001001100110011001100", "010100001011001100110011001100", "010100001101001100110011001100", "010100001111001100110011001100", 
"010100010001001100110011001100", "010100010011001100110011001100", "010100010101001100110011001100", "010100010111001100110011001100", 
"010100011001001100110011001100", "010100011011001100110011001100", "010100011101001100110011001100", "010100011111001100110011001100", 
"010100100001001100110011001100", "010100100011001100110011001100", "010100100101001100110011001100", "010100100111001100110011001100", 
"010100101001001100110011001100", "010100101011001100110011001100", "010100101101001100110011001100", "010100101111001100110011001100", 
"010100110001001100110011001100", "010100110011001100110011001100", "010100110101001100110011001100", "010100110111001100110011001100", 
"010100111001001100110011001100", "010100111011001100110011001100", "010100111101001100110011001100", "010100111111001100110011001100", 
"010101000001001100110011001100", "010101000011001100110011001100", "010101000101001100110011001100", "010101000111001100110011001100", 
"010101001001001100110011001100", "010101001011001100110011001100", "010101001101001100110011001100", "010101001111001100110011001100", 
"010101010001001100110011001100", "010101010011001100110011001100", "010101010101001100110011001100", "010101010111001100110011001100", 
"010101011001001100110011001100", "010101011011001100110011001100", "010101011101001100110011001100", "010101011111001100110011001100", 
"010101100001001100110011001100", "010101100011001100110011001100", "010101100101001100110011001100", "010101100111001100110011001100", 
"010101101001001100110011001100", "010101101011001100110011001100", "010101101101001100110011001100", "010101101111001100110011001100", 
"010101110001001100110011001100", "010101110011001100110011001100", "010101110101001100110011001100", "010101110111001100110011001100", 
"010101111001001100110011001100", "010101111011001100110011001100", "010101111101001100110011001100", "010101111111001100110011001100", 
"010110000001001100110011001100", "010110000011001100110011001100", "010110000101001100110011001100", "010110000111001100110011001100", 
"010110001001001100110011001100", "010110001011001100110011001100", "010110001101001100110011001100", "010110001111001100110011001100", 
"010110010001001100110011001100", "010110010011001100110011001100", "010110010101001100110011001100", "010110010111001100110011001100", 
"010110011001001100110011001100", "010110011011001100110011001100", "010110011101001100110011001100", "010110011111001100110011001100", 
"010110100001001100110011001100", "010110100011001100110011001100", "010110100101001100110011001100", "010110100111001100110011001100", 
"010110101001001100110011001100", "010110101011001100110011001100", "010110101101001100110011001100", "010110101111001100110011001100", 
"010110110001001100110011001100", "010110110011001100110011001100", "010110110101001100110011001100", "010110110111001100110011001100", 
"010110111001001100110011001100", "010110111011001100110011001100", "010110111101001100110011001100", "010110111111001100110011001100", 
"010111000001001100110011001100", "010111000011001100110011001100", "010111000101001100110011001100", "010111000111001100110011001100", 
"010111001001001100110011001100", "010111001011001100110011001100", "010111001101001100110011001100", "010111001111001100110011001100", 
"010111010001001100110011001100", "010111010011001100110011001100", "010111010101001100110011001100", "010111010111001100110011001100", 
"010111011001001100110011001100", "010111011011001100110011001100", "010111011101001100110011001100", "010111011111001100110011001100", 
"010111100001001100110011001100", "010111100011001100110011001100", "010111100101001100110011001100", "010111100111001100110011001100", 
"010111101001001100110011001100", "010111101011001100110011001100", "010111101101001100110011001100", "010111101111001100110011001100", 
"010111110001001100110011001100", "010111110011001100110011001100", "010111110101001100110011001100", "010111110111001100110011001100", 
"010111111001001100110011001100", "010111111011001100110011001100", "010111111101001100110011001100", "010111111111001100110011001100", 
"011000000001001100110011001100", "011000000011001100110011001100", "011000000101001100110011001100", "011000000111001100110011001100", 
"011000001001001100110011001100", "011000001011001100110011001100", "011000001101001100110011001100", "011000001111001100110011001100", 
"011000010001001100110011001100", "011000010011001100110011001100", "011000010101001100110011001100", "011000010111001100110011001100", 
"011000011001001100110011001100", "011000011011001100110011001100", "011000011101001100110011001100", "011000011111001100110011001100", 
"011000100001001100110011001100", "011000100011001100110011001100", "011000100101001100110011001100", "011000100111001100110011001100", 
"011000101001001100110011001100", "011000101011001100110011001100", "011000101101001100110011001100", "011000101111001100110011001100", 
"011000110001001100110011001100", "011000110011001100110011001100", "011000110101001100110011001100", "011000110111001100110011001100", 
"011000111001001100110011001100", "011000111011001100110011001100", "011000111101001100110011001100", "011000111111001100110011001100", 
"011001000001001100110011001100", "011001000011001100110011001100", "011001000101001100110011001100", "011001000111001100110011001100", 
"011001001001001100110011001100", "011001001011001100110011001100", "011001001101001100110011001100", "011001001111001100110011001100", 
"011001010001001100110011001100", "011001010011001100110011001100", "011001010101001100110011001100", "011001010111001100110011001100", 
"011001011001001100110011001100", "011001011011001100110011001100", "011001011101001100110011001100", "011001011111001100110011001100", 
"011001100001001100110011001100", "011001100011001100110011001100", "011001100101001100110011001100", "011001100111001100110011001100", 
"011001101001001100110011001100", "011001101011001100110011001100", "011001101101001100110011001100", "011001101111001100110011001100", 
"011001110001001100110011001100", "011001110011001100110011001100", "011001110101001100110011001100", "011001110111001100110011001100", 
"011001111001001100110011001100", "011001111011001100110011001100", "011001111101001100110011001100", "011001111111001100110011001100", 
"011010000001001100110011001100", "011010000011001100110011001100", "011010000101001100110011001100", "011010000111001100110011001100", 
"011010001001001100110011001100", "011010001011001100110011001100", "011010001101001100110011001100", "011010001111001100110011001100", 
"011010010001001100110011001100", "011010010011001100110011001100", "011010010101001100110011001100", "011010010111001100110011001100", 
"011010011001001100110011001100", "011010011011001100110011001100", "011010011101001100110011001100", "011010011111001100110011001100", 
"011010100001001100110011001100", "011010100011001100110011001100", "011010100101001100110011001100", "011010100111001100110011001100", 
"011010101001001100110011001100", "011010101011001100110011001100", "011010101101001100110011001100", "011010101111001100110011001100", 
"011010110001001100110011001100", "011010110011001100110011001100", "011010110101001100110011001100", "011010110111001100110011001100", 
"011010111001001100110011001100", "011010111011001100110011001100", "011010111101001100110011001100", "011010111111001100110011001100", 
"011011000001001100110011001100", "011011000011001100110011001100", "011011000101001100110011001100", "011011000111001100110011001100", 
"011011001001001100110011001100", "011011001011001100110011001100", "011011001101001100110011001100", "011011001111001100110011001100", 
"011011010001001100110011001100", "011011010011001100110011001100", "011011010101001100110011001100", "011011010111001100110011001100", 
"011011011001001100110011001100", "011011011011001100110011001100", "011011011101001100110011001100", "011011011111001100110011001100", 
"011011100001001100110011001100", "011011100011001100110011001100", "011011100101001100110011001100", "011011100111001100110011001100", 
"011011101001001100110011001100", "011011101011001100110011001100", "011011101101001100110011001100", "011011101111001100110011001100", 
"011011110001001100110011001100", "011011110011001100110011001100", "011011110101001100110011001100", "011011110111001100110011001100", 
"011011111001001100110011001100", "011011111011001100110011001100", "011011111101001100110011001100", "011011111111001100110011001100", 
"011100000001001100110011001100", "011100000011001100110011001100", "011100000101001100110011001100", "011100000111001100110011001100", 
"011100001001001100110011001100", "011100001011001100110011001100", "011100001101001100110011001100", "011100001111001100110011001100", 
"011100010001001100110011001100", "011100010011001100110011001100", "011100010101001100110011001100", "011100010111001100110011001100", 
"011100011001001100110011001100", "011100011011001100110011001100", "011100011101001100110011001100", "011100011111001100110011001100", 
"011100100001001100110011001100", "011100100011001100110011001100", "011100100101001100110011001100", "011100100111001100110011001100", 
"011100101001001100110011001100", "011100101011001100110011001100", "011100101101001100110011001100", "011100101111001100110011001100", 
"011100110001001100110011001100", "011100110011001100110011001100", "011100110101001100110011001100", "011100110111001100110011001100", 
"011100111001001100110011001100", "011100111011001100110011001100", "011100111101001100110011001100", "011100111111001100110011001100", 
"011101000001001100110011001100", "011101000011001100110011001100", "011101000101001100110011001100", "011101000111001100110011001100", 
"011101001001001100110011001100", "011101001011001100110011001100", "011101001101001100110011001100", "011101001111001100110011001100", 
"011101010001001100110011001100", "011101010011001100110011001100", "011101010101001100110011001100", "011101010111001100110011001100", 
"011101011001001100110011001100", "011101011011001100110011001100", "011101011101001100110011001100", "011101011111001100110011001100", 
"011101100001001100110011001100", "011101100011001100110011001100", "011101100101001100110011001100", "011101100111001100110011001100", 
"011101101001001100110011001100", "011101101011001100110011001100", "011101101101001100110011001100", "011101101111001100110011001100", 
"011101110001001100110011001100", "011101110011001100110011001100", "011101110101001100110011001100", "011101110111001100110011001100", 
"011101111001001100110011001100", "011101111011001100110011001100", "011101111101001100110011001100", "011101111111001100110011001100", 
"011110000001001100110011001100", "011110000011001100110011001100", "011110000101001100110011001100", "011110000111001100110011001100", 
"011110001001001100110011001100", "011110001011001100110011001100", "011110001101001100110011001100", "011110001111001100110011001100", 
"011110010001001100110011001100", "011110010011001100110011001100", "011110010101001100110011001100", "011110010111001100110011001100", 
"011110011001001100110011001100", "011110011011001100110011001100", "011110011101001100110011001100", "011110011111001100110011001100", 
"011110100001001100110011001100", "011110100011001100110011001100", "011110100101001100110011001100", "011110100111001100110011001100", 
"011110101001001100110011001100", "011110101011001100110011001100", "011110101101001100110011001100", "011110101111001100110011001100", 
"011110110001001100110011001100", "011110110011001100110011001100", "011110110101001100110011001100", "011110110111001100110011001100", 
"011110111001001100110011001100", "011110111011001100110011001100", "011110111101001100110011001100", "011110111111001100110011001100", 
"011111000001001100110011001100", "011111000011001100110011001100", "011111000101001100110011001100", "011111000111001100110011001100", 
"011111001001001100110011001100", "011111001011001100110011001100", "011111001101001100110011001100", "011111001111001100110011001100", 
"011111010001001100110011001100", "011111010011001100110011001100", "011111010101001100110011001100", "011111010111001100110011001100", 
"011111011001001100110011001100", "011111011011001100110011001100", "011111011101001100110011001100", "011111011111001100110011001100", 
"011111100001001100110011001100", "011111100011001100110011001100", "011111100101001100110011001100", "011111100111001100110011001100", 
"011111101001001100110011001100", "011111101011001100110011001100", "011111101101001100110011001100", "011111101111001100110011001100", 
"011111110001001100110011001100", "011111110011001100110011001100", "011111110101001100110011001100", "011111110111001100110011001100", 
"011111111001001100110011001100", "011111111011001100110011001100", "011111111101001100110011001100", "011111111111001100110011001100", 
"100000000001001100110011001100", "100000000011001100110011001100", "100000000101001100110011001100", "100000000111001100110011001100", 
"100000001001001100110011001100", "100000001011001100110011001100", "100000001101001100110011001100", "100000001111001100110011001100", 
"100000010001001100110011001100", "100000010011001100110011001100", "100000010101001100110011001100", "100000010111001100110011001100", 
"100000011001001100110011001100", "100000011011001100110011001100", "100000011101001100110011001100", "100000011111001100110011001100", 
"100000100001001100110011001100", "100000100011001100110011001100", "100000100101001100110011001100", "100000100111001100110011001100", 
"100000101001001100110011001100", "100000101011001100110011001100", "100000101101001100110011001100", "100000101111001100110011001100", 
"100000110001001100110011001100", "100000110011001100110011001100", "100000110101001100110011001100", "100000110111001100110011001100", 
"100000111001001100110011001100", "100000111011001100110011001100", "100000111101001100110011001100", "100000111111001100110011001100", 
"100001000001001100110011001100", "100001000011001100110011001100", "100001000101001100110011001100", "100001000111001100110011001100", 
"100001001001001100110011001100", "100001001011001100110011001100", "100001001101001100110011001100", "100001001111001100110011001100", 
"100001010001001100110011001100", "100001010011001100110011001100", "100001010101001100110011001100", "100001010111001100110011001100", 
"100001011001001100110011001100", "100001011011001100110011001100", "100001011101001100110011001100", "100001011111001100110011001100", 
"100001100001001100110011001100", "100001100011001100110011001100", "100001100101001100110011001100", "100001100111001100110011001100", 
"100001101001001100110011001100", "100001101011001100110011001100", "100001101101001100110011001100", "100001101111001100110011001100", 
"100001110001001100110011001100", "100001110011001100110011001100", "100001110101001100110011001100", "100001110111001100110011001100", 
"100001111001001100110011001100", "100001111011001100110011001100", "100001111101001100110011001100", "100001111111001100110011001100", 
"100010000001001100110011001100", "100010000011001100110011001100", "100010000101001100110011001100", "100010000111001100110011001100", 
"100010001001001100110011001100", "100010001011001100110011001100", "100010001101001100110011001100", "100010001111001100110011001100", 
"100010010001001100110011001100", "100010010011001100110011001100", "100010010101001100110011001100", "100010010111001100110011001100", 
"100010011001001100110011001100", "100010011011001100110011001100", "100010011101001100110011001100", "100010011111001100110011001100", 
"100010100001001100110011001100", "100010100011001100110011001100", "100010100101001100110011001100", "100010100111001100110011001100", 
"100010101001001100110011001100", "100010101011001100110011001100", "100010101101001100110011001100", "100010101111001100110011001100", 
"100010110001001100110011001100", "100010110011001100110011001100", "100010110101001100110011001100", "100010110111001100110011001100", 
"100010111001001100110011001100", "100010111011001100110011001100", "100010111101001100110011001100", "100010111111001100110011001100", 
"100011000001001100110011001100", "100011000011001100110011001100", "100011000101001100110011001100", "100011000111001100110011001100", 
"100011001001001100110011001100", "100011001011001100110011001100", "100011001101001100110011001100", "100011001111001100110011001100", 
"100011010001001100110011001100", "100011010011001100110011001100", "100011010101001100110011001100", "100011010111001100110011001100", 
"100011011001001100110011001100", "100011011011001100110011001100", "100011011101001100110011001100", "100011011111001100110011001100", 
"100011100001001100110011001100", "100011100011001100110011001100", "100011100101001100110011001100", "100011100111001100110011001100", 
"100011101001001100110011001100", "100011101011001100110011001100", "100011101101001100110011001100", "100011101111001100110011001100", 
"100011110001001100110011001100", "100011110011001100110011001100", "100011110101001100110011001100", "100011110111001100110011001100", 
"100011111001001100110011001100", "100011111011001100110011001100", "100011111101001100110011001100", "100011111111001100110011001100", 
"100100000001001100110011001100", "100100000011001100110011001100", "100100000101001100110011001100", "100100000111001100110011001100", 
"100100001001001100110011001100", "100100001011001100110011001100", "100100001101001100110011001100", "100100001111001100110011001100", 
"100100010001001100110011001100", "100100010011001100110011001100", "100100010101001100110011001100", "100100010111001100110011001100", 
"100100011001001100110011001100", "100100011011001100110011001100", "100100011101001100110011001100", "100100011111001100110011001100", 
"100100100001001100110011001100", "100100100011001100110011001100", "100100100101001100110011001100", "100100100111001100110011001100", 
"100100101001001100110011001100", "100100101011001100110011001100", "100100101101001100110011001100", "100100101111001100110011001100", 
"100100110001001100110011001100", "100100110011001100110011001100", "100100110101001100110011001100", "100100110111001100110011001100", 
"100100111001001100110011001100", "100100111011001100110011001100", "100100111101001100110011001100", "100100111111001100110011001100", 
"100101000001001100110011001100", "100101000011001100110011001100", "100101000101001100110011001100", "100101000111001100110011001100", 
"100101001001001100110011001100", "100101001011001100110011001100", "100101001101001100110011001100", "100101001111001100110011001100", 
"100101010001001100110011001100", "100101010011001100110011001100", "100101010101001100110011001100", "100101010111001100110011001100", 
"100101011001001100110011001100", "100101011011001100110011001100", "100101011101001100110011001100", "100101011111001100110011001100", 
"100101100001001100110011001100", "100101100011001100110011001100", "100101100101001100110011001100", "100101100111001100110011001100", 
"100101101001001100110011001100", "100101101011001100110011001100", "100101101101001100110011001100", "100101101111001100110011001100", 
"100101110001001100110011001100", "100101110011001100110011001100", "100101110101001100110011001100", "100101110111001100110011001100", 
"100101111001001100110011001100", "100101111011001100110011001100", "100101111101001100110011001100", "100101111111001100110011001100", 
"100110000001001100110011001100", "100110000011001100110011001100", "100110000101001100110011001100", "100110000111001100110011001100", 
"100110001001001100110011001100", "100110001011001100110011001100", "100110001101001100110011001100", "100110001111001100110011001100", 
"100110010001001100110011001100", "100110010011001100110011001100", "100110010101001100110011001100", "100110010111001100110011001100", 
"100110011001001100110011001100", "100110011011001100110011001100", "100110011101001100110011001100", "100110011111001100110011001100", 
"100110100001001100110011001100", "100110100011001100110011001100", "100110100101001100110011001100", "100110100111001100110011001100", 
"100110101001001100110011001100", "100110101011001100110011001100", "100110101101001100110011001100", "100110101111001100110011001100", 
"100110110001001100110011001100", "100110110011001100110011001100", "100110110101001100110011001100", "100110110111001100110011001100", 
"100110111001001100110011001100", "100110111011001100110011001100", "100110111101001100110011001100", "100110111111001100110011001100", 
"100111000001001100110011001100", "100111000011001100110011001100", "100111000101001100110011001100", "100111000111001100110011001100", 
"100111001001001100110011001100", "100111001011001100110011001100", "100111001101001100110011001100", "100111001111001100110011001100", 
"100111010001001100110011001100", "100111010011001100110011001100", "100111010101001100110011001100", "100111010111001100110011001100", 
"100111011001001100110011001100", "100111011011001100110011001100", "100111011101001100110011001100", "100111011111001100110011001100", 
"100111100001001100110011001100", "100111100011001100110011001100", "100111100101001100110011001100", "100111100111001100110011001100", 
"100111101001001100110011001100", "100111101011001100110011001100", "100111101101001100110011001100", "100111101111001100110011001100", 
"100111110001001100110011001100", "100111110011001100110011001100", "100111110101001100110011001100", "100111110111001100110011001100", 
"100111111001001100110011001100", "100111111011001100110011001100", "100111111101001100110011001100", "100111111111001100110011001100", 
"101000000001001100110011001100", "101000000011001100110011001100", "101000000101001100110011001100", "101000000111001100110011001100", 
"101000001001001100110011001100", "101000001011001100110011001100", "101000001101001100110011001100", "101000001111001100110011001100", 
"101000010001001100110011001100", "101000010011001100110011001100", "101000010101001100110011001100", "101000010111001100110011001100", 
"101000011001001100110011001100", "101000011011001100110011001100", "101000011101001100110011001100", "101000011111001100110011001100", 
"101000100001001100110011001100", "101000100011001100110011001100", "101000100101001100110011001100", "101000100111001100110011001100", 
"101000101001001100110011001100", "101000101011001100110011001100", "101000101101001100110011001100", "101000101111001100110011001100", 
"101000110001001100110011001100", "101000110011001100110011001100", "101000110101001100110011001100", "101000110111001100110011001100", 
"101000111001001100110011001100", "101000111011001100110011001100", "101000111101001100110011001100", "101000111111001100110011001100", 
"101001000001001100110011001100", "101001000011001100110011001100", "101001000101001100110011001100", "101001000111001100110011001100", 
"101001001001001100110011001100", "101001001011001100110011001100", "101001001101001100110011001100", "101001001111001100110011001100", 
"101001010001001100110011001100", "101001010011001100110011001100", "101001010101001100110011001100", "101001010111001100110011001100", 
"101001011001001100110011001100", "101001011011001100110011001100", "101001011101001100110011001100", "101001011111001100110011001100", 
"101001100001001100110011001100", "101001100011001100110011001100", "101001100101001100110011001100", "101001100111001100110011001100", 
"101001101001001100110011001100", "101001101011001100110011001100", "101001101101001100110011001100", "101001101111001100110011001100", 
"101001110001001100110011001100", "101001110011001100110011001100", "101001110101001100110011001100", "101001110111001100110011001100", 
"101001111001001100110011001100", "101001111011001100110011001100", "101001111101001100110011001100", "101001111111001100110011001100", 
"101010000001001100110011001100", "101010000011001100110011001100", "101010000101001100110011001100", "101010000111001100110011001100", 
"101010001001001100110011001100", "101010001011001100110011001100", "101010001101001100110011001100", "101010001111001100110011001100", 
"101010010001001100110011001100", "101010010011001100110011001100", "101010010101001100110011001100", "101010010111001100110011001100", 
"101010011001001100110011001100", "101010011011001100110011001100", "101010011101001100110011001100", "101010011111001100110011001100", 
"101010100001001100110011001100", "101010100011001100110011001100", "101010100101001100110011001100", "101010100111001100110011001100", 
"101010101001001100110011001100", "101010101011001100110011001100", "101010101101001100110011001100", "101010101111001100110011001100", 
"101010110001001100110011001100", "101010110011001100110011001100", "101010110101001100110011001100", "101010110111001100110011001100", 
"101010111001001100110011001100", "101010111011001100110011001100", "101010111101001100110011001100", "101010111111001100110011001100", 
"101011000001001100110011001100", "101011000011001100110011001100", "101011000101001100110011001100", "101011000111001100110011001100", 
"101011001001001100110011001100", "101011001011001100110011001100", "101011001101001100110011001100", "101011001111001100110011001100", 
"101011010001001100110011001100", "101011010011001100110011001100", "101011010101001100110011001100", "101011010111001100110011001100", 
"101011011001001100110011001100", "101011011011001100110011001100", "101011011101001100110011001100", "101011011111001100110011001100", 
"101011100001001100110011001100", "101011100011001100110011001100", "101011100101001100110011001100", "101011100111001100110011001100", 
"101011101001001100110011001100", "101011101011001100110011001100", "101011101101001100110011001100", "101011101111001100110011001100", 
"101011110001001100110011001100", "101011110011001100110011001100", "101011110101001100110011001100", "101011110111001100110011001100", 
"101011111001001100110011001100", "101011111011001100110011001100", "101011111101001100110011001100", "101011111111001100110011001100", 
"101100000001001100110011001100", "101100000011001100110011001100", "101100000101001100110011001100", "101100000111001100110011001100", 
"101100001001001100110011001100", "101100001011001100110011001100", "101100001101001100110011001100", "101100001111001100110011001100", 
"101100010001001100110011001100", "101100010011001100110011001100", "101100010101001100110011001100", "101100010111001100110011001100", 
"101100011001001100110011001100", "101100011011001100110011001100", "101100011101001100110011001100", "101100011111001100110011001100", 
"101100100001001100110011001100", "101100100011001100110011001100", "101100100101001100110011001100", "101100100111001100110011001100", 
"101100101001001100110011001100", "101100101011001100110011001100", "101100101101001100110011001100", "101100101111001100110011001100", 
"101100110001001100110011001100", "101100110011001100110011001100", "101100110101001100110011001100", "101100110111001100110011001100", 
"101100111001001100110011001100", "101100111011001100110011001100", "101100111101001100110011001100", "101100111111001100110011001100", 
"101101000001001100110011001100", "101101000011001100110011001100", "101101000101001100110011001100", "101101000111001100110011001100", 
"101101001001001100110011001100", "101101001011001100110011001100", "101101001101001100110011001100", "101101001111001100110011001100", 
"101101010001001100110011001100", "101101010011001100110011001100", "101101010101001100110011001100", "101101010111001100110011001100", 
"101101011001001100110011001100", "101101011011001100110011001100", "101101011101001100110011001100", "101101011111001100110011001100", 
"101101100001001100110011001100", "101101100011001100110011001100", "101101100101001100110011001100", "101101100111001100110011001100", 
"101101101001001100110011001100", "101101101011001100110011001100", "101101101101001100110011001100", "101101101111001100110011001100", 
"101101110001001100110011001100", "101101110011001100110011001100", "101101110101001100110011001100", "101101110111001100110011001100", 
"101101111001001100110011001100", "101101111011001100110011001100", "101101111101001100110011001100", "101101111111001100110011001100", 
"101110000001001100110011001100", "101110000011001100110011001100", "101110000101001100110011001100", "101110000111001100110011001100", 
"101110001001001100110011001100", "101110001011001100110011001100", "101110001101001100110011001100", "101110001111001100110011001100", 
"101110010001001100110011001100", "101110010011001100110011001100", "101110010101001100110011001100", "101110010111001100110011001100", 
"101110011001001100110011001100", "101110011011001100110011001100", "101110011101001100110011001100", "101110011111001100110011001100", 
"101110100001001100110011001100", "101110100011001100110011001100", "101110100101001100110011001100", "101110100111001100110011001100", 
"101110101001001100110011001100", "101110101011001100110011001100", "101110101101001100110011001100", "101110101111001100110011001100", 
"101110110001001100110011001100", "101110110011001100110011001100", "101110110101001100110011001100", "101110110111001100110011001100", 
"101110111001001100110011001100", "101110111011001100110011001100", "101110111101001100110011001100", "101110111111001100110011001100", 
"101111000001001100110011001100", "101111000011001100110011001100", "101111000101001100110011001100", "101111000111001100110011001100", 
"101111001001001100110011001100", "101111001011001100110011001100", "101111001101001100110011001100", "101111001111001100110011001100", 
"101111010001001100110011001100", "101111010011001100110011001100", "101111010101001100110011001100", "101111010111001100110011001100", 
"101111011001001100110011001100", "101111011011001100110011001100", "101111011101001100110011001100", "101111011111001100110011001100", 
"101111100001001100110011001100", "101111100011001100110011001100", "101111100101001100110011001100", "101111100111001100110011001100", 
"101111101001001100110011001100", "101111101011001100110011001100", "101111101101001100110011001100", "101111101111001100110011001100", 
"101111110001001100110011001100", "101111110011001100110011001100", "101111110101001100110011001100", "101111110111001100110011001100", 
"101111111001001100110011001100", "101111111011001100110011001100", "101111111101001100110011001100", "101111111111001100110011001100", 
"110000000001001100110011001100", "110000000011001100110011001100", "110000000101001100110011001100", "110000000111001100110011001100", 
"110000001001001100110011001100", "110000001011001100110011001100", "110000001101001100110011001100", "110000001111001100110011001100", 
"110000010001001100110011001100", "110000010011001100110011001100", "110000010101001100110011001100", "110000010111001100110011001100", 
"110000011001001100110011001100", "110000011011001100110011001100", "110000011101001100110011001100", "110000011111001100110011001100", 
"110000100001001100110011001100", "110000100011001100110011001100", "110000100101001100110011001100", "110000100111001100110011001100", 
"110000101001001100110011001100", "110000101011001100110011001100", "110000101101001100110011001100", "110000101111001100110011001100", 
"110000110001001100110011001100", "110000110011001100110011001100", "110000110101001100110011001100", "110000110111001100110011001100", 
"110000111001001100110011001100", "110000111011001100110011001100", "110000111101001100110011001100", "110000111111001100110011001100", 
"110001000001001100110011001100", "110001000011001100110011001100", "110001000101001100110011001100", "110001000111001100110011001100", 
"110001001001001100110011001100", "110001001011001100110011001100", "110001001101001100110011001100", "110001001111001100110011001100", 
"110001010001001100110011001100", "110001010011001100110011001100", "110001010101001100110011001100", "110001010111001100110011001100", 
"110001011001001100110011001100", "110001011011001100110011001100", "110001011101001100110011001100", "110001011111001100110011001100", 
"110001100001001100110011001100", "110001100011001100110011001100", "110001100101001100110011001100", "110001100111001100110011001100", 
"110001101001001100110011001100", "110001101011001100110011001100", "110001101101001100110011001100", "110001101111001100110011001100", 
"110001110001001100110011001100", "110001110011001100110011001100", "110001110101001100110011001100", "110001110111001100110011001100", 
"110001111001001100110011001100", "110001111011001100110011001100", "110001111101001100110011001100", "110001111111001100110011001100", 
"110010000001001100110011001100", "110010000011001100110011001100", "110010000101001100110011001100", "110010000111001100110011001100", 
"110010001001001100110011001100", "110010001011001100110011001100", "110010001101001100110011001100", "110010001111001100110011001100", 
"110010010001001100110011001100", "110010010011001100110011001100", "110010010101001100110011001100", "110010010111001100110011001100", 
"110010011001001100110011001100", "110010011011001100110011001100", "110010011101001100110011001100", "110010011111001100110011001100", 
"110010100001001100110011001100", "110010100011001100110011001100", "110010100101001100110011001100", "110010100111001100110011001100", 
"110010101001001100110011001100", "110010101011001100110011001100", "110010101101001100110011001100", "110010101111001100110011001100", 
"110010110001001100110011001100", "110010110011001100110011001100", "110010110101001100110011001100", "110010110111001100110011001100", 
"110010111001001100110011001100", "110010111011001100110011001100", "110010111101001100110011001100", "110010111111001100110011001100", 
"110011000001001100110011001100", "110011000011001100110011001100", "110011000101001100110011001100", "110011000111001100110011001100", 
"110011001001001100110011001100", "110011001011001100110011001100", "110011001101001100110011001100", "110011001111001100110011001100", 
"110011010001001100110011001100", "110011010011001100110011001100", "110011010101001100110011001100", "110011010111001100110011001100", 
"110011011001001100110011001100", "110011011011001100110011001100", "110011011101001100110011001100", "110011011111001100110011001100", 
"110011100001001100110011001100", "110011100011001100110011001100", "110011100101001100110011001100", "110011100111001100110011001100", 
"110011101001001100110011001100", "110011101011001100110011001100", "110011101101001100110011001100", "110011101111001100110011001100", 
"110011110001001100110011001100", "110011110011001100110011001100", "110011110101001100110011001100", "110011110111001100110011001100", 
"110011111001001100110011001100", "110011111011001100110011001100", "110011111101001100110011001100", "110011111111001100110011001100", 
"110100000001001100110011001100", "110100000011001100110011001100", "110100000101001100110011001100", "110100000111001100110011001100", 
"110100001001001100110011001100", "110100001011001100110011001100", "110100001101001100110011001100", "110100001111001100110011001100", 
"110100010001001100110011001100", "110100010011001100110011001100", "110100010101001100110011001100", "110100010111001100110011001100", 
"110100011001001100110011001100", "110100011011001100110011001100", "110100011101001100110011001100", "110100011111001100110011001100", 
"110100100001001100110011001100", "110100100011001100110011001100", "110100100101001100110011001100", "110100100111001100110011001100", 
"110100101001001100110011001100", "110100101011001100110011001100", "110100101101001100110011001100", "110100101111001100110011001100", 
"110100110001001100110011001100", "110100110011001100110011001100", "110100110101001100110011001100", "110100110111001100110011001100", 
"110100111001001100110011001100", "110100111011001100110011001100", "110100111101001100110011001100", "110100111111001100110011001100", 
"110101000001001100110011001100", "110101000011001100110011001100", "110101000101001100110011001100", "110101000111001100110011001100", 
"110101001001001100110011001100", "110101001011001100110011001100", "110101001101001100110011001100", "110101001111001100110011001100", 
"110101010001001100110011001100", "110101010011001100110011001100", "110101010101001100110011001100", "110101010111001100110011001100", 
"110101011001001100110011001100", "110101011011001100110011001100", "110101011101001100110011001100", "110101011111001100110011001100", 
"110101100001001100110011001100", "110101100011001100110011001100", "110101100101001100110011001100", "110101100111001100110011001100", 
"110101101001001100110011001100", "110101101011001100110011001100", "110101101101001100110011001100", "110101101111001100110011001100", 
"110101110001001100110011001100", "110101110011001100110011001100", "110101110101001100110011001100", "110101110111001100110011001100", 
"110101111001001100110011001100", "110101111011001100110011001100", "110101111101001100110011001100", "110101111111001100110011001100", 
"110110000001001100110011001100", "110110000011001100110011001100", "110110000101001100110011001100", "110110000111001100110011001100", 
"110110001001001100110011001100", "110110001011001100110011001100", "110110001101001100110011001100", "110110001111001100110011001100", 
"110110010001001100110011001100", "110110010011001100110011001100", "110110010101001100110011001100", "110110010111001100110011001100", 
"110110011001001100110011001100", "110110011011001100110011001100", "110110011101001100110011001100", "110110011111001100110011001100", 
"110110100001001100110011001100", "110110100011001100110011001100", "110110100101001100110011001100", "110110100111001100110011001100", 
"110110101001001100110011001100", "110110101011001100110011001100", "110110101101001100110011001100", "110110101111001100110011001100", 
"110110110001001100110011001100", "110110110011001100110011001100", "110110110101001100110011001100", "110110110111001100110011001100", 
"110110111001001100110011001100", "110110111011001100110011001100", "110110111101001100110011001100", "110110111111001100110011001100", 
"110111000001001100110011001100", "110111000011001100110011001100", "110111000101001100110011001100", "110111000111001100110011001100", 
"110111001001001100110011001100", "110111001011001100110011001100", "110111001101001100110011001100", "110111001111001100110011001100", 
"110111010001001100110011001100", "110111010011001100110011001100", "110111010101001100110011001100", "110111010111001100110011001100", 
"110111011001001100110011001100", "110111011011001100110011001100", "110111011101001100110011001100", "110111011111001100110011001100", 
"110111100001001100110011001100", "110111100011001100110011001100", "110111100101001100110011001100", "110111100111001100110011001100", 
"110111101001001100110011001100", "110111101011001100110011001100", "110111101101001100110011001100", "110111101111001100110011001100", 
"110111110001001100110011001100", "110111110011001100110011001100", "110111110101001100110011001100", "110111110111001100110011001100", 
"110111111001001100110011001100", "110111111011001100110011001100", "110111111101001100110011001100", "110111111111001100110011001100", 
"111000000001001100110011001100", "111000000011001100110011001100", "111000000101001100110011001100", "111000000111001100110011001100", 
"111000001001001100110011001100", "111000001011001100110011001100", "111000001101001100110011001100", "111000001111001100110011001100", 
"111000010001001100110011001100", "111000010011001100110011001100", "111000010101001100110011001100", "111000010111001100110011001100", 
"111000011001001100110011001100", "111000011011001100110011001100", "111000011101001100110011001100", "111000011111001100110011001100", 
"111000100001001100110011001100", "111000100011001100110011001100", "111000100101001100110011001100", "111000100111001100110011001100", 
"111000101001001100110011001100", "111000101011001100110011001100", "111000101101001100110011001100", "111000101111001100110011001100", 
"111000110001001100110011001100", "111000110011001100110011001100", "111000110101001100110011001100", "111000110111001100110011001100", 
"111000111001001100110011001100", "111000111011001100110011001100", "111000111101001100110011001100", "111000111111001100110011001100", 
"111001000001001100110011001100", "111001000011001100110011001100", "111001000101001100110011001100", "111001000111001100110011001100", 
"111001001001001100110011001100", "111001001011001100110011001100", "111001001101001100110011001100", "111001001111001100110011001100", 
"111001010001001100110011001100", "111001010011001100110011001100", "111001010101001100110011001100", "111001010111001100110011001100", 
"111001011001001100110011001100", "111001011011001100110011001100", "111001011101001100110011001100", "111001011111001100110011001100", 
"111001100001001100110011001100", "111001100011001100110011001100", "111001100101001100110011001100", "111001100111001100110011001100", 
"111001101001001100110011001100", "111001101011001100110011001100", "111001101101001100110011001100", "111001101111001100110011001100", 
"111001110001001100110011001100", "111001110011001100110011001100", "111001110101001100110011001100", "111001110111001100110011001100", 
"111001111001001100110011001100", "111001111011001100110011001100", "111001111101001100110011001100", "111001111111001100110011001100", 
"111010000001001100110011001100", "111010000011001100110011001100", "111010000101001100110011001100", "111010000111001100110011001100", 
"111010001001001100110011001100", "111010001011001100110011001100", "111010001101001100110011001100", "111010001111001100110011001100", 
"111010010001001100110011001100", "111010010011001100110011001100", "111010010101001100110011001100", "111010010111001100110011001100", 
"111010011001001100110011001100", "111010011011001100110011001100", "111010011101001100110011001100", "111010011111001100110011001100", 
"111010100001001100110011001100", "111010100011001100110011001100", "111010100101001100110011001100", "111010100111001100110011001100", 
"111010101001001100110011001100", "111010101011001100110011001100", "111010101101001100110011001100", "111010101111001100110011001100", 
"111010110001001100110011001100", "111010110011001100110011001100", "111010110101001100110011001100", "111010110111001100110011001100", 
"111010111001001100110011001100", "111010111011001100110011001100", "111010111101001100110011001100", "111010111111001100110011001100", 
"111011000001001100110011001100", "111011000011001100110011001100", "111011000101001100110011001100", "111011000111001100110011001100", 
"111011001001001100110011001100", "111011001011001100110011001100", "111011001101001100110011001100", "111011001111001100110011001100", 
"111011010001001100110011001100", "111011010011001100110011001100", "111011010101001100110011001100", "111011010111001100110011001100", 
"111011011001001100110011001100", "111011011011001100110011001100", "111011011101001100110011001100", "111011011111001100110011001100", 
"111011100001001100110011001100", "111011100011001100110011001100", "111011100101001100110011001100", "111011100111001100110011001100", 
"111011101001001100110011001100", "111011101011001100110011001100", "111011101101001100110011001100", "111011101111001100110011001100", 
"111011110001001100110011001100", "111011110011001100110011001100", "111011110101001100110011001100", "111011110111001100110011001100", 
"111011111001001100110011001100", "111011111011001100110011001100", "111011111101001100110011001100", "111011111111001100110011001100", 
"111100000001001100110011001100", "111100000011001100110011001100", "111100000101001100110011001100", "111100000111001100110011001100", 
"111100001001001100110011001100", "111100001011001100110011001100", "111100001101001100110011001100", "111100001111001100110011001100", 
"111100010001001100110011001100", "111100010011001100110011001100", "111100010101001100110011001100", "111100010111001100110011001100", 
"111100011001001100110011001100", "111100011011001100110011001100", "111100011101001100110011001100", "111100011111001100110011001100", 
"111100100001001100110011001100", "111100100011001100110011001100", "111100100101001100110011001100", "111100100111001100110011001100", 
"111100101001001100110011001100", "111100101011001100110011001100", "111100101101001100110011001100", "111100101111001100110011001100", 
"111100110001001100110011001100", "111100110011001100110011001100", "111100110101001100110011001100", "111100110111001100110011001100", 
"111100111001001100110011001100", "111100111011001100110011001100", "111100111101001100110011001100", "111100111111001100110011001100", 
"111101000001001100110011001100", "111101000011001100110011001100", "111101000101001100110011001100", "111101000111001100110011001100", 
"111101001001001100110011001100", "111101001011001100110011001100", "111101001101001100110011001100", "111101001111001100110011001100", 
"111101010001001100110011001100", "111101010011001100110011001100", "111101010101001100110011001100", "111101010111001100110011001100", 
"111101011001001100110011001100", "111101011011001100110011001100", "111101011101001100110011001100", "111101011111001100110011001100", 
"111101100001001100110011001100", "111101100011001100110011001100", "111101100101001100110011001100", "111101100111001100110011001100", 
"111101101001001100110011001100", "111101101011001100110011001100", "111101101101001100110011001100", "111101101111001100110011001100", 
"111101110001001100110011001100", "111101110011001100110011001100", "111101110101001100110011001100", "111101110111001100110011001100", 
"111101111001001100110011001100", "111101111011001100110011001100", "111101111101001100110011001100", "111101111111001100110011001100", 
"111110000001001100110011001100", "111110000011001100110011001100", "111110000101001100110011001100", "111110000111001100110011001100", 
"111110001001001100110011001100", "111110001011001100110011001100", "111110001101001100110011001100", "111110001111001100110011001100", 
"111110010001001100110011001100", "111110010011001100110011001100", "111110010101001100110011001100", "111110010111001100110011001100", 
"111110011001001100110011001100", "111110011011001100110011001100", "111110011101001100110011001100", "111110011111001100110011001100", 
"111110100001001100110011001100", "111110100011001100110011001100", "111110100101001100110011001100", "111110100111001100110011001100", 
"111110101001001100110011001100", "111110101011001100110011001100", "111110101101001100110011001100", "111110101111001100110011001100", 
"111110110001001100110011001100", "111110110011001100110011001100", "111110110101001100110011001100", "111110110111001100110011001100", 
"111110111001001100110011001100", "111110111011001100110011001100", "111110111101001100110011001100", "111110111111001100110011001100", 
"111111000001001100110011001100", "111111000011001100110011001100", "111111000101001100110011001100", "111111000111001100110011001100", 
"111111001001001100110011001100", "111111001011001100110011001100", "111111001101001100110011001100", "111111001111001100110011001100", 
"111111010001001100110011001100", "111111010011001100110011001100", "111111010101001100110011001100", "111111010111001100110011001100", 
"111111011001001100110011001100", "111111011011001100110011001100", "111111011101001100110011001100", "111111011111001100110011001100", 
"111111100001001100110011001100", "111111100011001100110011001100", "111111100101001100110011001100", "111111100111001100110011001100", 
"111111101001001100110011001100", "111111101011001100110011001100", "111111101101001100110011001100", "111111101111001100110011001100", 
"111111110001001100110011001100", "111111110011001100110011001100", "111111110101001100110011001100", "111111110111001100110011001100", 
"111111111001001100110011001100", "111111111011001100110011001100", "111111111101001100110011001100", "111111111111001100110011001100"
);
type muon_pt_lut_ufixed_array is array (0 to 2**(D_S_I_MUON_V2.pt_high-D_S_I_MUON_V2.pt_low+1)-1) of ufixed(7 downto -20);
constant MU_PT_LUT_UFIXED : muon_pt_lut_ufixed_array := (
"0000000000000000000000000000", "0000000001001100110011001100", "0000000011001100110011001100", "0000000101001100110011001100", 
"0000000111001100110011001100", "0000001001001100110011001100", "0000001011001100110011001100", "0000001101001100110011001100", 
"0000001111001100110011001100", "0000010001001100110011001100", "0000010011001100110011001100", "0000010101001100110011001100", 
"0000010111001100110011001100", "0000011001001100110011001100", "0000011011001100110011001100", "0000011101001100110011001100", 
"0000011111001100110011001100", "0000100001001100110011001100", "0000100011001100110011001100", "0000100101001100110011001100", 
"0000100111001100110011001100", "0000101001001100110011001100", "0000101011001100110011001100", "0000101101001100110011001100", 
"0000101111001100110011001100", "0000110001001100110011001100", "0000110011001100110011001100", "0000110101001100110011001100", 
"0000110111001100110011001100", "0000111001001100110011001100", "0000111011001100110011001100", "0000111101001100110011001100", 
"0000111111001100110011001100", "0001000001001100110011001100", "0001000011001100110011001100", "0001000101001100110011001100", 
"0001000111001100110011001100", "0001001001001100110011001100", "0001001011001100110011001100", "0001001101001100110011001100", 
"0001001111001100110011001100", "0001010001001100110011001100", "0001010011001100110011001100", "0001010101001100110011001100", 
"0001010111001100110011001100", "0001011001001100110011001100", "0001011011001100110011001100", "0001011101001100110011001100", 
"0001011111001100110011001100", "0001100001001100110011001100", "0001100011001100110011001100", "0001100101001100110011001100", 
"0001100111001100110011001100", "0001101001001100110011001100", "0001101011001100110011001100", "0001101101001100110011001100", 
"0001101111001100110011001100", "0001110001001100110011001100", "0001110011001100110011001100", "0001110101001100110011001100", 
"0001110111001100110011001100", "0001111001001100110011001100", "0001111011001100110011001100", "0001111101001100110011001100", 
"0001111111001100110011001100", "0010000001001100110011001100", "0010000011001100110011001100", "0010000101001100110011001100", 
"0010000111001100110011001100", "0010001001001100110011001100", "0010001011001100110011001100", "0010001101001100110011001100", 
"0010001111001100110011001100", "0010010001001100110011001100", "0010010011001100110011001100", "0010010101001100110011001100", 
"0010010111001100110011001100", "0010011001001100110011001100", "0010011011001100110011001100", "0010011101001100110011001100", 
"0010011111001100110011001100", "0010100001001100110011001100", "0010100011001100110011001100", "0010100101001100110011001100", 
"0010100111001100110011001100", "0010101001001100110011001100", "0010101011001100110011001100", "0010101101001100110011001100", 
"0010101111001100110011001100", "0010110001001100110011001100", "0010110011001100110011001100", "0010110101001100110011001100", 
"0010110111001100110011001100", "0010111001001100110011001100", "0010111011001100110011001100", "0010111101001100110011001100", 
"0010111111001100110011001100", "0011000001001100110011001100", "0011000011001100110011001100", "0011000101001100110011001100", 
"0011000111001100110011001100", "0011001001001100110011001100", "0011001011001100110011001100", "0011001101001100110011001100", 
"0011001111001100110011001100", "0011010001001100110011001100", "0011010011001100110011001100", "0011010101001100110011001100", 
"0011010111001100110011001100", "0011011001001100110011001100", "0011011011001100110011001100", "0011011101001100110011001100", 
"0011011111001100110011001100", "0011100001001100110011001100", "0011100011001100110011001100", "0011100101001100110011001100", 
"0011100111001100110011001100", "0011101001001100110011001100", "0011101011001100110011001100", "0011101101001100110011001100", 
"0011101111001100110011001100", "0011110001001100110011001100", "0011110011001100110011001100", "0011110101001100110011001100", 
"0011110111001100110011001100", "0011111001001100110011001100", "0011111011001100110011001100", "0011111101001100110011001100", 
"0011111111001100110011001100", "0100000001001100110011001100", "0100000011001100110011001100", "0100000101001100110011001100", 
"0100000111001100110011001100", "0100001001001100110011001100", "0100001011001100110011001100", "0100001101001100110011001100", 
"0100001111001100110011001100", "0100010001001100110011001100", "0100010011001100110011001100", "0100010101001100110011001100", 
"0100010111001100110011001100", "0100011001001100110011001100", "0100011011001100110011001100", "0100011101001100110011001100", 
"0100011111001100110011001100", "0100100001001100110011001100", "0100100011001100110011001100", "0100100101001100110011001100", 
"0100100111001100110011001100", "0100101001001100110011001100", "0100101011001100110011001100", "0100101101001100110011001100", 
"0100101111001100110011001100", "0100110001001100110011001100", "0100110011001100110011001100", "0100110101001100110011001100", 
"0100110111001100110011001100", "0100111001001100110011001100", "0100111011001100110011001100", "0100111101001100110011001100", 
"0100111111001100110011001100", "0101000001001100110011001100", "0101000011001100110011001100", "0101000101001100110011001100", 
"0101000111001100110011001100", "0101001001001100110011001100", "0101001011001100110011001100", "0101001101001100110011001100", 
"0101001111001100110011001100", "0101010001001100110011001100", "0101010011001100110011001100", "0101010101001100110011001100", 
"0101010111001100110011001100", "0101011001001100110011001100", "0101011011001100110011001100", "0101011101001100110011001100", 
"0101011111001100110011001100", "0101100001001100110011001100", "0101100011001100110011001100", "0101100101001100110011001100", 
"0101100111001100110011001100", "0101101001001100110011001100", "0101101011001100110011001100", "0101101101001100110011001100", 
"0101101111001100110011001100", "0101110001001100110011001100", "0101110011001100110011001100", "0101110101001100110011001100", 
"0101110111001100110011001100", "0101111001001100110011001100", "0101111011001100110011001100", "0101111101001100110011001100", 
"0101111111001100110011001100", "0110000001001100110011001100", "0110000011001100110011001100", "0110000101001100110011001100", 
"0110000111001100110011001100", "0110001001001100110011001100", "0110001011001100110011001100", "0110001101001100110011001100", 
"0110001111001100110011001100", "0110010001001100110011001100", "0110010011001100110011001100", "0110010101001100110011001100", 
"0110010111001100110011001100", "0110011001001100110011001100", "0110011011001100110011001100", "0110011101001100110011001100", 
"0110011111001100110011001100", "0110100001001100110011001100", "0110100011001100110011001100", "0110100101001100110011001100", 
"0110100111001100110011001100", "0110101001001100110011001100", "0110101011001100110011001100", "0110101101001100110011001100", 
"0110101111001100110011001100", "0110110001001100110011001100", "0110110011001100110011001100", "0110110101001100110011001100", 
"0110110111001100110011001100", "0110111001001100110011001100", "0110111011001100110011001100", "0110111101001100110011001100", 
"0110111111001100110011001100", "0111000001001100110011001100", "0111000011001100110011001100", "0111000101001100110011001100", 
"0111000111001100110011001100", "0111001001001100110011001100", "0111001011001100110011001100", "0111001101001100110011001100", 
"0111001111001100110011001100", "0111010001001100110011001100", "0111010011001100110011001100", "0111010101001100110011001100", 
"0111010111001100110011001100", "0111011001001100110011001100", "0111011011001100110011001100", "0111011101001100110011001100", 
"0111011111001100110011001100", "0111100001001100110011001100", "0111100011001100110011001100", "0111100101001100110011001100", 
"0111100111001100110011001100", "0111101001001100110011001100", "0111101011001100110011001100", "0111101101001100110011001100", 
"0111101111001100110011001100", "0111110001001100110011001100", "0111110011001100110011001100", "0111110101001100110011001100", 
"0111110111001100110011001100", "0111111001001100110011001100", "0111111011001100110011001100", "0111111101001100110011001100", 
"0111111111001100110011001100", "1000000001001100110011001100", "1000000011001100110011001100", "1000000101001100110011001100", 
"1000000111001100110011001100", "1000001001001100110011001100", "1000001011001100110011001100", "1000001101001100110011001100", 
"1000001111001100110011001100", "1000010001001100110011001100", "1000010011001100110011001100", "1000010101001100110011001100", 
"1000010111001100110011001100", "1000011001001100110011001100", "1000011011001100110011001100", "1000011101001100110011001100", 
"1000011111001100110011001100", "1000100001001100110011001100", "1000100011001100110011001100", "1000100101001100110011001100", 
"1000100111001100110011001100", "1000101001001100110011001100", "1000101011001100110011001100", "1000101101001100110011001100", 
"1000101111001100110011001100", "1000110001001100110011001100", "1000110011001100110011001100", "1000110101001100110011001100", 
"1000110111001100110011001100", "1000111001001100110011001100", "1000111011001100110011001100", "1000111101001100110011001100", 
"1000111111001100110011001100", "1001000001001100110011001100", "1001000011001100110011001100", "1001000101001100110011001100", 
"1001000111001100110011001100", "1001001001001100110011001100", "1001001011001100110011001100", "1001001101001100110011001100", 
"1001001111001100110011001100", "1001010001001100110011001100", "1001010011001100110011001100", "1001010101001100110011001100", 
"1001010111001100110011001100", "1001011001001100110011001100", "1001011011001100110011001100", "1001011101001100110011001100", 
"1001011111001100110011001100", "1001100001001100110011001100", "1001100011001100110011001100", "1001100101001100110011001100", 
"1001100111001100110011001100", "1001101001001100110011001100", "1001101011001100110011001100", "1001101101001100110011001100", 
"1001101111001100110011001100", "1001110001001100110011001100", "1001110011001100110011001100", "1001110101001100110011001100", 
"1001110111001100110011001100", "1001111001001100110011001100", "1001111011001100110011001100", "1001111101001100110011001100", 
"1001111111001100110011001100", "1010000001001100110011001100", "1010000011001100110011001100", "1010000101001100110011001100", 
"1010000111001100110011001100", "1010001001001100110011001100", "1010001011001100110011001100", "1010001101001100110011001100", 
"1010001111001100110011001100", "1010010001001100110011001100", "1010010011001100110011001100", "1010010101001100110011001100", 
"1010010111001100110011001100", "1010011001001100110011001100", "1010011011001100110011001100", "1010011101001100110011001100", 
"1010011111001100110011001100", "1010100001001100110011001100", "1010100011001100110011001100", "1010100101001100110011001100", 
"1010100111001100110011001100", "1010101001001100110011001100", "1010101011001100110011001100", "1010101101001100110011001100", 
"1010101111001100110011001100", "1010110001001100110011001100", "1010110011001100110011001100", "1010110101001100110011001100", 
"1010110111001100110011001100", "1010111001001100110011001100", "1010111011001100110011001100", "1010111101001100110011001100", 
"1010111111001100110011001100", "1011000001001100110011001100", "1011000011001100110011001100", "1011000101001100110011001100", 
"1011000111001100110011001100", "1011001001001100110011001100", "1011001011001100110011001100", "1011001101001100110011001100", 
"1011001111001100110011001100", "1011010001001100110011001100", "1011010011001100110011001100", "1011010101001100110011001100", 
"1011010111001100110011001100", "1011011001001100110011001100", "1011011011001100110011001100", "1011011101001100110011001100", 
"1011011111001100110011001100", "1011100001001100110011001100", "1011100011001100110011001100", "1011100101001100110011001100", 
"1011100111001100110011001100", "1011101001001100110011001100", "1011101011001100110011001100", "1011101101001100110011001100", 
"1011101111001100110011001100", "1011110001001100110011001100", "1011110011001100110011001100", "1011110101001100110011001100", 
"1011110111001100110011001100", "1011111001001100110011001100", "1011111011001100110011001100", "1011111101001100110011001100", 
"1011111111001100110011001100", "1100000001001100110011001100", "1100000011001100110011001100", "1100000101001100110011001100", 
"1100000111001100110011001100", "1100001001001100110011001100", "1100001011001100110011001100", "1100001101001100110011001100", 
"1100001111001100110011001100", "1100010001001100110011001100", "1100010011001100110011001100", "1100010101001100110011001100", 
"1100010111001100110011001100", "1100011001001100110011001100", "1100011011001100110011001100", "1100011101001100110011001100", 
"1100011111001100110011001100", "1100100001001100110011001100", "1100100011001100110011001100", "1100100101001100110011001100", 
"1100100111001100110011001100", "1100101001001100110011001100", "1100101011001100110011001100", "1100101101001100110011001100", 
"1100101111001100110011001100", "1100110001001100110011001100", "1100110011001100110011001100", "1100110101001100110011001100", 
"1100110111001100110011001100", "1100111001001100110011001100", "1100111011001100110011001100", "1100111101001100110011001100", 
"1100111111001100110011001100", "1101000001001100110011001100", "1101000011001100110011001100", "1101000101001100110011001100", 
"1101000111001100110011001100", "1101001001001100110011001100", "1101001011001100110011001100", "1101001101001100110011001100", 
"1101001111001100110011001100", "1101010001001100110011001100", "1101010011001100110011001100", "1101010101001100110011001100", 
"1101010111001100110011001100", "1101011001001100110011001100", "1101011011001100110011001100", "1101011101001100110011001100", 
"1101011111001100110011001100", "1101100001001100110011001100", "1101100011001100110011001100", "1101100101001100110011001100", 
"1101100111001100110011001100", "1101101001001100110011001100", "1101101011001100110011001100", "1101101101001100110011001100", 
"1101101111001100110011001100", "1101110001001100110011001100", "1101110011001100110011001100", "1101110101001100110011001100", 
"1101110111001100110011001100", "1101111001001100110011001100", "1101111011001100110011001100", "1101111101001100110011001100", 
"1101111111001100110011001100", "1110000001001100110011001100", "1110000011001100110011001100", "1110000101001100110011001100", 
"1110000111001100110011001100", "1110001001001100110011001100", "1110001011001100110011001100", "1110001101001100110011001100", 
"1110001111001100110011001100", "1110010001001100110011001100", "1110010011001100110011001100", "1110010101001100110011001100", 
"1110010111001100110011001100", "1110011001001100110011001100", "1110011011001100110011001100", "1110011101001100110011001100", 
"1110011111001100110011001100", "1110100001001100110011001100", "1110100011001100110011001100", "1110100101001100110011001100", 
"1110100111001100110011001100", "1110101001001100110011001100", "1110101011001100110011001100", "1110101101001100110011001100", 
"1110101111001100110011001100", "1110110001001100110011001100", "1110110011001100110011001100", "1110110101001100110011001100", 
"1110110111001100110011001100", "1110111001001100110011001100", "1110111011001100110011001100", "1110111101001100110011001100", 
"1110111111001100110011001100", "1111000001001100110011001100", "1111000011001100110011001100", "1111000101001100110011001100", 
"1111000111001100110011001100", "1111001001001100110011001100", "1111001011001100110011001100", "1111001101001100110011001100", 
"1111001111001100110011001100", "1111010001001100110011001100", "1111010011001100110011001100", "1111010101001100110011001100", 
"1111010111001100110011001100", "1111011001001100110011001100", "1111011011001100110011001100", "1111011101001100110011001100", 
"1111011111001100110011001100", "1111100001001100110011001100", "1111100011001100110011001100", "1111100101001100110011001100", 
"1111100111001100110011001100", "1111101001001100110011001100", "1111101011001100110011001100", "1111101101001100110011001100", 
"1111101111001100110011001100", "1111110001001100110011001100", "1111110011001100110011001100", "1111110101001100110011001100", 
"1111110111001100110011001100", "1111111001001100110011001100", "1111111011001100110011001100", "1111111101001100110011001100"
);
type calo_calo_diff_eta_lut_ufixed_array is array (0 to 2**MAX_CALO_ETA_BITS-1) of ufixed(3 downto -20);
constant CALO_CALO_DIFF_ETA_LUT_UFIXED : calo_calo_diff_eta_lut_ufixed_array := (
"000000000000000000000000", "000000001011010000111000", "000000010110010001011010", "000000100001100010010010", 
"000000101100100010110100", "000000110111100011010100", "000001000010110100001110", "000001001110000101000110", 
"000001011001000101101000", "000001100100000110001000", "000001101111010111000010", "000001111010100111111010", 
"000010000101101000011100", "000010010000111001010110", "000010011011111001110110", "000010100111001010110000", 
"000010110010001011010000", "000010111101001011110000", "000011001000011100101010", "000011010011011101001010", 
"000011011110101110000100", "000011101001111110111110", "000011110100111111011110", "000100000000010000011000", 
"000100001011010000111000", "000100010110100001110010", "000100100001100010010010", "000100101100100010110100", 
"000100110111110011101100", "000101000010110100001110", "000101001110000101000110", "000101011001000101101000", 
"000101100100010110100000", "000101101111100111011010", "000101111010100111111010", "000110000101111000110100", 
"000110010000111001010110", "000110011100001010001110", "000110100111001010110000", "000110110010011011101000", 
"000110111101011100001010", "000111001000011100101010", "000111010011101101100100", "000111011110101110000100", 
"000111101001111110111110", "000111110100111111011110", "001000000000010000011000", "001000001011010000111000", 
"001000010110100001110010", "001000100001110010101100", "001000101100110011001100", "001000110111110011101100", 
"001001000011000100100110", "001001001110010101100000", "001001011001010110000000", "001001100100010110100000", 
"001001101111100111011010", "001001111010111000010100", "001010000101111000110100", "001010010001001001101110", 
"001010011100001010001110", "001010100111001010110000", "001010110010011011101000", "001010111101101100100010", 
"001011001000101101000010", "001011010011101101100100", "001011011110111110011100", "001011101010001111010110", 
"001011110101001111110110", "001100000000010000011000", "001100001011100001010000", "001100010110110010001010", 
"001100100001110010101100", "001100101101000011100100", "001100111000000100000110", "001101000011000100100110", 
"001101001110010101100000", "001101011001100110011000", "001101100100100110111010", "001101101111100111011010", 
"001101111010111000010100", "001110000110001001001100", "001110010001001001101110", "001110011100001010001110", 
"001110100111011011001000", "001110110010101100000010", "001110111101101100100010", "001111001000101101000010", 
"001111010011111101111100", "001111011110111110011100", "001111101010001111010110", "001111110101100000010000", 
"010000000000100000110000", "010000001011100001010000", "010000010110110010001010", "010000100001110010101100", 
"010000101101000011100100", "010000111000010100011110", "010001000011010100111110", "010001001110100101111000", 
"010001011001100110011000", "010001100100100110111010", "010001101111110111110010", "010001111010111000010100", 
"010010000110001001001100", "010010010001011010000110", "010010011100011010100110", "010010100111101011100000", 
"010010110010101100000010", "010010111101101100100010", "010011001000111101011100", "010011010100001110010100", 
"010011011111001110110110", "010011101010011111101110", "010011110101100000010000", "010100000000100000110000", 
"010100001011110001101010", "010100010110110010001010", "010100100010000011000100", "010100101101010011111100", 
"010100111000010100011110", "010101000011100101011000", "010101001110100101111000", "010101011001100110011000", 
"010101100100110111010010", "010101110000001000001100", "010101111011001000101100", "010110000110011001100110", 
"010110010001011010000110", "010110011100011010100110", "010110100111101011100000", "010110110010101100000010", 
"010110111101111100111010", "010111001001001101110100", "010111010100001110010100", "010111011111011111001110", 
"010111101010011111101110", "010111110101100000010000", "011000000000110001001000", "011000001100000010000010", 
"011000010111000010100010", "011000100010010011011100", "011000101101010011111100", "011000111000010100011110", 
"011001000011100101011000", "011001001110100101111000", "011001011001110110110010", "011001100101000111101010", 
"011001110000001000001100", "011001111011011001000100", "011010000110011001100110", "011010010001011010000110", 
"011010011100101011000000", "011010100111111011111000", "011010110010111100011010", "011010111110001101010010", 
"011011001001001101110100", "011011010100001110010100", "011011011111011111001110", "011011101010011111101110", 
"011011110101110000101000", "011100000001000001100010", "011100001100000010000010", "011100010111010010111100", 
"011100100010010011011100", "011100101101010011111100", "011100111000100100110110", "011101000011100101011000", 
"011101001110110110010000", "011101011010000111001010", "011101100101000111101010", "011101110000001000001100", 
"011101111011011001000100", "011110000110011001100110", "011110010001101010011110", "011110011100111011011000", 
"011110100111111011111000", "011110110011001100110010", "011110111110001101010010", "011111001001001101110100", 
"011111010100011110101110", "011111011111011111001110", "011111101010110000001000", "011111110110000001000000", 
"100000000001000001100010", "100000001100000010000010", "100000010111010010111100", "100000100010010011011100", 
"100000101101100100010110", "100000111000100100110110", "100001000011110101110000", "100001001110110110010000", 
"100001011010000111001010", "100001100101011000000100", "100001110000011000100100", "100001111011101001011110", 
"100010000110101001111110", "100010010001111010111000", "100010011100111011011000", "100010101000001100010010", 
"100010110011001100110010", "100010111110011101101100", "100011001001011110001100", "100011010100011110101110", 
"100011011111101111100110", "100011101010110000001000", "100011110110000001000000", "100100000001010001111010", 
"100100001100010010011010", "100100010111100011010100", "100100100010100011110100", "100100101101110100101110", 
"100100111000110101001110", "100101000100000110001000", "100101001111000110101000", "100101011010010111100010", 
"100101100101011000000100", "100101110000011000100100", "100101111011101001011110", "100110000110101001111110", 
"100110010001111010111000", "100110011101001011110000", "100110101000001100010010", "100110110011011101001010", 
"100110111110011101101100", "100111001001101110100100", "100111010100101111000110", "100111011111111111111110", 
"100111101011000000100000", "100111110110010001011010", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000"
);
type calo_calo_diff_phi_lut_ufixed_array is array (0 to 2**MAX_CALO_PHI_BITS-1) of ufixed(2 downto -20);
constant CALO_CALO_DIFF_PHI_LUT_UFIXED : calo_calo_diff_phi_lut_ufixed_array := (
"00000000000000000000000", "00000001011010000111000", "00000010110010001011010", "00000100001100010010010", 
"00000101100110011001100", "00000110111110011101100", "00001000011000100100110", "00001001110000101000110", 
"00001011001010110000000", "00001100100100110111010", "00001101111100111011010", "00001111010111000010100", 
"00010000110001001001100", "00010010001001001101110", "00010011100011010100110", "00010100111011011001000", 
"00010110010101100000010", "00010111101111100111010", "00011001000111101011100", "00011010100001110010100", 
"00011011111011111001110", "00011101010011111101110", "00011110101110000101000", "00100000001000001100010", 
"00100001100000010000010", "00100010111010010111100", "00100100010010011011100", "00100101101100100010110", 
"00100111000110101001110", "00101000011110101110000", "00101001111000110101000", "00101011010010111100010", 
"00101100101011000000100", "00101110000101000111100", "00101111011111001110110", "00110000110111010010110", 
"00110010010001011010000", "00110011101001011110000", "00110101000011100101010", "00110110011101101100100", 
"00110111110101110000100", "00111001001111110111110", "00111010101001111110110", "00111100000010000011000", 
"00111101011100001010000", "00111110110100001110010", "01000000001110010101100", "01000001101000011100100", 
"01000011000000100000110", "01000100011010100111110", "01000101110100101111000", "01000111001100110011000", 
"01001000100110111010010", "01001010000001000001100", "01001011011001000101100", "01001100110011001100110", 
"01001110001011010000110", "01001111100101011000000", "01010000111111011111000", "01010010010111100011010", 
"01010011110001101010010", "01010101001011110001100", "01010110100011110101110", "01010111111101111100110", 
"01011001011000000100000", "01011010110000001000000", "01011100001010001111010", "01011101100010010011010", 
"01011110111100011010100", "01100000010110100001110", "01100001101110100101110", "01100011001000101101000", 
"01100100100010110100000", "01100101111010111000010", "01100111010100111111010", "01101000101101000011100", 
"01101010000111001010110", "01101011100001010001110", "01101100111001010110000", "01101110010011011101000", 
"01101111101101100100010", "01110001000101101000010", "01110010011111101111100", "01110011111001110110110", 
"01110101010001111010110", "01110110101100000010000", "01111000000100000110000", "01111001011110001101010", 
"01111010111000010100010", "01111100010000011000100", "01111101101010011111100", "01111111000100100110110", 
"10000000011100101011000", "10000001110110110010000", "10000011010000111001010", "10000100101000111101010", 
"10000110000011000100100", "10000111011011001000100", "10001000110101001111110", "10001010001111010111000", 
"10001011100111011011000", "10001101000001100010010", "10001110011011101001010", "10001111110011101101100", 
"10010001001101110100100", "10010010100101111000110", "10010011111111111111110", "10010101011010000111000", 
"10010110110010001011010", "10011000001100010010010", "10011001100110011001100", "10011010111110011101100", 
"10011100011000100100110", "10011101110010101100000", "10011111001010110000000", "10100000100100110111010", 
"10100001111100111011010", "10100011010111000010100", "10100100110001001001100", "10100110001001001101110", 
"10100111100011010100110", "10101000111101011100000", "10101010010101100000010", "10101011101111100111010", 
"10101101001001101110100", "10101110100001110010100", "10101111111011111001110", "10110001010011111101110", 
"10110010101110000101000", "10110100001000001100010", "10110101100000010000010", "10110110111010010111100", 
"10111000010100011110100", "10111001101100100010110", "10111011000110101001110", "10111100011110101110000", 
"10111101111000110101000", "10111111010010111100010", "11000000101011000000100", "11000010000101000111100", 
"11000011011111001110110", "11000100110111010010110", "11000110010001011010000", "11000111101011100001010", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000"
);
type calo_calo_cosh_deta_lut_ufixed_array is array (0 to 2**MAX_CALO_ETA_BITS-1) of ufixed(13 downto -20);
constant CALO_CALO_COSH_DETA_LUT_UFIXED : calo_calo_cosh_deta_lut_ufixed_array := (
"0000000000000100000000000000000000", "0000000000000100000000010000011000", "0000000000000100000001000001100010", "0000000000000100000010010011011100", 
"0000000000000100000011110101110000", "0000000000000100000110001001001100", "0000000000000100001000101101000010", "0000000000000100001100000010000010", 
"0000000000000100001111100111011010", "0000000000000100010011111101111100", "0000000000000100011000100100110110", "0000000000000100011101111100111010", 
"0000000000000100100011100101011000", "0000000000000100101001111110111110", "0000000000000100110000111001010110", "0000000000000100111000100100110110", 
"0000000000000101000000100000110000", "0000000000000101001001001101110100", "0000000000000101010010101100000010", "0000000000000101011100011010100110", 
"0000000000000101100111001010110000", "0000000000000101110010011011101000", "0000000000000101111110011101101100", "0000000000000110001011010000111000", 
"0000000000000110011000100100110110", "0000000000000110100110111010010110", "0000000000000110110110000001000000", "0000000000000111000101111000110100", 
"0000000000000111010110100001110010", "0000000000000111101000001100010010", "0000000000000111111010100111111010", "0000000000001000001110010101100000", 
"0000000000001000100010110100001110", "0000000000001000111000010100011110", "0000000000001001001110110110010000", "0000000000001001100110101001111110", 
"0000000000001001111111011111001110", "0000000000001010011001100110011000", "0000000000001010110100111111011110", "0000000000001011010001101010011110", 
"0000000000001011101111100111011010", "0000000000001100001111000110101000", "0000000000001100110000001000001100", "0000000000001101010010101100000010", 
"0000000000001101110110110010001010", "0000000000001110011100011010100110", "0000000000001111000100000110001000", "0000000000001111101101010011111100", 
"0000000000010000011000100100110110", "0000000000010001000101111000110100", "0000000000010001110101001111110110", "0000000000010010100110101001111110", 
"0000000000010011011010010111100010", "0000000000010100010000011000100100", "0000000000010101001000111101011100", "0000000000010110000100000110001000", 
"0000000000010111000001110010101100", "0000000000011000000010100011110100", "0000000000011001000101111000110100", "0000000000011010001100010010011010", 
"0000000000011011010110000001000000", "0000000000011100100011000100100110", "0000000000011101110011011101001010", "0000000000011111000111101011100000", 
"0000000000100000011111011111001110", "0000000000100001111011001000101100", "0000000000100011011011001000101100", "0000000000100100111111001110110110", 
"0000000000100110100111111011111000", "0000000000101000010101001111110110", "0000000000101010000111011011001000", "0000000000101011111110101110000100", 
"0000000000101101111011011001000100", "0000000000101111111101011100001010", "0000000000110010000101101000011100", "0000000000110100010011101101100100", 
"0000000000110110100111111011111000", "0000000000111001000011000100100110", "0000000000111011100100110111010010", "0000000000111110001110000101000110", 
"0000000001000000111110101110000100", "0000000001000011110111010010111100", "0000000001000110111000000100000110", "0000000001001010000001100010010010", 
"0000000001001101010011101101100100", "0000000001010000101111100111011010", "0000000001010100010100111111011110", "0000000001011000000100100110111010", 
"0000000001011011111110111110011100", "0000000001100000000100100110111010", "0000000001100100010101110000101000", "0000000001101000110010111100011010", 
"0000000001101101011100111011011000", "0000000001110010010100001110010100", "0000000001110111011001000101101000", "0000000001111100101100110011001100", 
"0000000010000010001111010111000010", "0000000010001000000001110010101100", "0000000010001110000100100110111010", "0000000010010100011000110101001110", 
"0000000010011010111110111110011100", "0000000010100001110111110011101100", "0000000010101001000100000110001000", "0000000010110000100101000111101010", 
"0000000010111000011011011001000100", "0000000011000000101000001100010010", "0000000011001001001100000010000010", "0000000011010010001000011100101010", 
"0000000011011011011110001101010010", "0000000011100101001110100101111000", "0000000011101111011010111000010100", "0000000011111010000100000110001000", 
"0000000100000101001011100001010000", "0000000100010000110010011011101000", "0000000100011100111010100111111010", "0000000100101001100101011000000100", 
"0000000100110110110011111101111100", "0000000101000100101000001100010010", "0000000101010011000011110101110000", "0000000101100010001000101101000010", 
"0000000101110001111000010100011110", "0000000110000010010100101111000110", "0000000110010011011111111111111110", "0000000110100101011011111001110110", 
"0000000110111000001011000000100000", "0000000111001011101111100111011010", "0000000111100000001011100001010000", "0000000111110101100001110010101100", 
"0000001000001011110100111111011110", "0000001000100011000111011011001000", "0000001000111011011100001010001110", "0000001001010100110110000001000000", 
"0000001001101111011000010100011110", "0000001010001011000110001001001100", "0000001010101000000010110100001110", "0000001011000110010001101010011110", 
"0000001011100101110110110010001010", "0000001100000110110101100000010000", "0000001100101001010010011011101000", "0000001101001101010001001001101110", 
"0000001101110010110110010001011010", "0000001110011010000110011001100110", "0000001111000011000110001001001100", "0000001111101101111010010111100010", 
"0000010000011010101000101101000010", "0000010001001001010110010001011010", "0000010001111010001000101101000010", "0000010010101101000101111000110100", 
"0000010011100010010011111101111100", "0000010100011001111001110110110010", "0000010101010011111101101100100010", "0000010110010000100110101001111110", 
"0000010111001111111100001010001110", "0000011000010010000110001001001100", "0000011001010111001100010010011010", "0000011010011111010110110010001010", 
"0000011011101010101110110110010000", "0000011100111001011101011100001010", "0000011110001011101011110001101010", "0000011111100001100100010110100000", 
"0000100000111011010001001001101110", "0000100010011000111101011100001010", "0000100011111010110011111101111100", "0000100101100001000001000001100010", 
"0000100111001011110001001001101110", "0000101000111011010000101000111100", "0000101010101111101101100100010110", "0000101100101001010110000001000000", 
"0000101110101000011000010100011110", "0000110000101101000100010110100000", "0000110010110111101001101110100100", "0000110101001000011001010110000000", 
"0000110111011111100101000111101010", "0000111001111101011110101110000100", "0000111100100010011001110110110010", "0000111111001110101010001111010110", 
"0001000010000010100100110111010010", "0001000100111110011111001110110110", "0001001000000010110000011000100100", "0001001011001111110000001000001100", 
"0001001110100101110111000010100010", "0001010010000101011111001110110110", "0001010101101111000011100101011000", "0001011001100011000000110001001000", 
"0001011101100001110011111101111100", "0001100001101011111100001010001110", "0001100110000001111001110110110010", "0001101010100100001110000101000110", 
"0001101111010011011100101011000000", "0001110100010000001001111110111110", "0001111001011010111100101011000000", "0001111110110100011100011010100110", 
"0010000100011101010011001100110010", "0010001010010110001100110011001100", "0010010000011111110110110010001010", "0010010110111011000001000001100010", 
"0010011101101000011101001011110000", "0010100100101000111111011111001110", "0010101011111101011101101100100010", "0010110011100110110001001001101110", 
"0010111011100101110100101111000110", "0011000011111011100110101001111110", "0011001100101001000111011011001000", "0011010101101111011010010111100010", 
"0011011111001111100110011001100110", "0011101001001010110100101111000110", "0011110011100010010010101100000010", "0011111110010111010000101000111100", 
"0100001001101011000010010011011100", "0100010101011110111111011111001110", "0100100001110100100011100101011000", "0100101110101101001110010101100000", 
"0100111100001010100011100101011000", "0101001010001110001011110001101010", "0101011000111001110011111101111100", "0101101000001111001101100100010110", 
"0101111000010000001111110111110010", "0110001000111110110110110010001010", "0110011010011101000100000110001000", "0110101100101100111110111110011100", 
"0110111111110000110101001111110110", "0111010011101010111010100111111010", "0111101000011101101001001101110100", "0111111110001011100010010011011100", 
"1000010100110111001110010101100000", "1000101100100011011100111011011000", "1001000101010011000101111000110100", "1001011111001001001001001101110100", 
"1001111010001000101110110110010000", "1010010110010101001000001100010010", "0000000000000000000000000000000000", "0000000000000000000000000000000000", 
"0000000000000000000000000000000000", "0000000000000000000000000000000000", "0000000000000000000000000000000000", "0000000000000000000000000000000000", 
"0000000000000000000000000000000000", "0000000000000000000000000000000000", "0000000000000000000000000000000000", "0000000000000000000000000000000000", 
"0000000000000000000000000000000000", "0000000000000000000000000000000000", "0000000000000000000000000000000000", "0000000000000000000000000000000000", 
"0000000000000000000000000000000000", "0000000000000000000000000000000000", "0000000000000000000000000000000000", "0000000000000000000000000000000000", 
"0000000000000000000000000000000000", "0000000000000000000000000000000000", "0000000000000000000000000000000000", "0000000000000000000000000000000000", 
"0000000000000000000000000000000000", "0000000000000000000000000000000000", "0000000000000000000000000000000000", "0000000000000000000000000000000000"
);
type calo_calo_cos_dphi_lut_ufixed_array is array (0 to 2**MAX_CALO_PHI_BITS-1) of ufixed(0 downto -20);
constant CALO_CALO_COS_DPHI_LUT_UFIXED : calo_calo_cos_dphi_lut_ufixed_array := (
"100000000000000000000", "011111111101111100110", "011111110111110011100", "011111101101100100010", 
"011111100001010001110", "011111001110110110010", "011110111010010111100", "011110100001110010100", 
"011110000101000111100", "011101100100010110100", "011100111111011111000", "011100011000100100110", 
"011011101101100100010", "011010111110011101100", "011010001101010011110", "011001011000000100000", 
"011000100000110001000", "010111100101011000000", "010110100111111011110", "010101101000011100100", 
"010100100100110111010", "010011011111001110110", "010010010111100011010", "010001001011110001100", 
"001111111111111111110", "001110110010001011010", "001101100010010011010", "001100010000011000100", 
"001010111100011010100", "001001101000011100100", "001000010010011011100", "000110111010010111100", 
"000101100100010110100", "000100001100010010010", "000010110010001011010", "000001011010000111000", 
"000000000000000000000", "000001011010000111000", "000010110010001011010", "000100001100010010010", 
"000101100100010110100", "000110111010010111100", "001000010010011011100", "001001101000011100100", 
"001010111100011010100", "001100010000011000100", "001101100010010011010", "001110110010001011010", 
"001111111111111111110", "010001001011110001100", "010010010111100011010", "010011011111001110110", 
"010100100100110111010", "010101101000011100100", "010110100111111011110", "010111100101011000000", 
"011000100000110001000", "011001011000000100000", "011010001101010011110", "011010111110011101100", 
"011011101101100100010", "011100011000100100110", "011100111111011111000", "011101100100010110100", 
"011110000101000111100", "011110100001110010100", "011110111010010111100", "011111001110110110010", 
"011111100001010001110", "011111101101100100010", "011111110111110011100", "011111111101111100110", 
"100000000000000000000", "011111111101111100110", "011111110111110011100", "011111101101100100010", 
"011111100001010001110", "011111001110110110010", "011110111010010111100", "011110100001110010100", 
"011110000101000111100", "011101100100010110100", "011100111111011111000", "011100011000100100110", 
"011011101101100100010", "011010111110011101100", "011010001101010011110", "011001011000000100000", 
"011000100000110001000", "010111100101011000000", "010110100111111011110", "010101101000011100100", 
"010100100100110111010", "010011011111001110110", "010010010111100011010", "010001001011110001100", 
"001111111111111111110", "001110110010001011010", "001101100010010011010", "001100010000011000100", 
"001010111100011010100", "001001101000011100100", "001000010010011011100", "000110111010010111100", 
"000101100100010110100", "000100001100010010010", "000010110010001011010", "000001011010000111000", 
"000000000000000000000", "000001011010000111000", "000010110010001011010", "000100001100010010010", 
"000101100100010110100", "000110111010010111100", "001000010010011011100", "001001101000011100100", 
"001010111100011010100", "001100010000011000100", "001101100010010011010", "001110110010001011010", 
"001111111111111111110", "010001001011110001100", "010010010111100011010", "010011011111001110110", 
"010100100100110111010", "010101101000011100100", "010110100111111011110", "010111100101011000000", 
"011000100000110001000", "011001011000000100000", "011010001101010011110", "011010111110011101100", 
"011011101101100100010", "011100011000100100110", "011100111111011111000", "011101100100010110100", 
"011110000101000111100", "011110100001110010100", "011110111010010111100", "011111001110110110010", 
"011111100001010001110", "011111101101100100010", "011111110111110011100", "011111111101111100110", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000"
);
type calo_calo_cos_dphi_sign_lut_array is array (0 to 2**MAX_CALO_PHI_BITS-1) of boolean;
constant CALO_CALO_COS_DPHI_SIGN_LUT : calo_calo_cos_dphi_sign_lut_array := (
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false
);
type muon_muon_diff_eta_lut_ufixed_array is array (0 to 2**(MUON_ETA_HIGH-MUON_ETA_LOW+1)-1) of ufixed(2 downto -20);
constant MU_MU_DIFF_ETA_LUT_UFIXED : muon_muon_diff_eta_lut_ufixed_array := (
"00000000000000000000000", "00000000010110100001110", "00000000101101000011100", "00000001000011100101010", 
"00000001011010000111000", "00000001101110100101110", "00000010000101000111100", "00000010011011101001010", 
"00000010110010001011010", "00000011001000101101000", "00000011011111001110110", "00000011110101110000100", 
"00000100001100010010010", "00000100100000110001000", "00000100110111010010110", "00000101001101110100100", 
"00000101100100010110100", "00000101111010111000010", "00000110010001011010000", "00000110100111111011110", 
"00000110111100011010100", "00000111010010111100010", "00000111101001011110000", "00000111111111111111110", 
"00001000010110100001110", "00001000101101000011100", "00001001000011100101010", "00001001011010000111000", 
"00001001110000101000110", "00001010000101000111100", "00001010011011101001010", "00001010110010001011010", 
"00001011001000101101000", "00001011011111001110110", "00001011110101110000100", "00001100001100010010010", 
"00001100100000110001000", "00001100110111010010110", "00001101001101110100100", "00001101100100010110100", 
"00001101111010111000010", "00001110010001011010000", "00001110100111111011110", "00001110111110011101100", 
"00001111010100111111010", "00001111101001011110000", "00001111111111111111110", "00010000010110100001110", 
"00010000101101000011100", "00010001000011100101010", "00010001011010000111000", "00010001110000101000110", 
"00010010000111001010110", "00010010011011101001010", "00010010110010001011010", "00010011001000101101000", 
"00010011011111001110110", "00010011110101110000100", "00010100001100010010010", "00010100100010110100000", 
"00010100111001010110000", "00010101001101110100100", "00010101100100010110100", "00010101111010111000010", 
"00010110010001011010000", "00010110100111111011110", "00010110111110011101100", "00010111010100111111010", 
"00010111101001011110000", "00010111111111111111110", "00011000010110100001110", "00011000101101000011100", 
"00011001000011100101010", "00011001011010000111000", "00011001110000101000110", "00011010000111001010110", 
"00011010011011101001010", "00011010110010001011010", "00011011001000101101000", "00011011011111001110110", 
"00011011110101110000100", "00011100001100010010010", "00011100100010110100000", "00011100111001010110000", 
"00011101001111110111110", "00011101100100010110100", "00011101111010111000010", "00011110010001011010000", 
"00011110100111111011110", "00011110111110011101100", "00011111010100111111010", "00011111101011100001010", 
"00100000000010000011000", "00100000010110100001110", "00100000101101000011100", "00100001000011100101010", 
"00100001011010000111000", "00100001110000101000110", "00100010000111001010110", "00100010011101101100100", 
"00100010110100001110010", "00100011001000101101000", "00100011011111001110110", "00100011110101110000100", 
"00100100001100010010010", "00100100100010110100000", "00100100111001010110000", "00100101001111110111110", 
"00100101100100010110100", "00100101111010111000010", "00100110010001011010000", "00100110100111111011110", 
"00100110111110011101100", "00100111010100111111010", "00100111101011100001010", "00101000000010000011000", 
"00101000010110100001110", "00101000101101000011100", "00101001000011100101010", "00101001011010000111000", 
"00101001110000101000110", "00101010000111001010110", "00101010011101101100100", "00101010110100001110010", 
"00101011001000101101000", "00101011011111001110110", "00101011110101110000100", "00101100001100010010010", 
"00101100100010110100000", "00101100111001010110000", "00101101001111110111110", "00101101100110011001100", 
"00101101111100111011010", "00101110010001011010000", "00101110100111111011110", "00101110111110011101100", 
"00101111010100111111010", "00101111101011100001010", "00110000000010000011000", "00110000011000100100110", 
"00110000101111000110100", "00110001000011100101010", "00110001011010000111000", "00110001110000101000110", 
"00110010000111001010110", "00110010011101101100100", "00110010110100001110010", "00110011001010110000000", 
"00110011100001010001110", "00110011110101110000100", "00110100001100010010010", "00110100100010110100000", 
"00110100111001010110000", "00110101001111110111110", "00110101100110011001100", "00110101111100111011010", 
"00110110010011011101000", "00110110100111111011110", "00110110111110011101100", "00110111010100111111010", 
"00110111101011100001010", "00111000000010000011000", "00111000011000100100110", "00111000101111000110100", 
"00111001000011100101010", "00111001011010000111000", "00111001110000101000110", "00111010000111001010110", 
"00111010011101101100100", "00111010110100001110010", "00111011001010110000000", "00111011100001010001110", 
"00111011110101110000100", "00111100001100010010010", "00111100100010110100000", "00111100111001010110000", 
"00111101001111110111110", "00111101100110011001100", "00111101111100111011010", "00111110010011011101000", 
"00111110100111111011110", "00111110111110011101100", "00111111010100111111010", "00111111101011100001010", 
"01000000000010000011000", "01000000011000100100110", "01000000101111000110100", "01000001000101101000010", 
"01000001011010000111000", "01000001110000101000110", "01000010000111001010110", "01000010011101101100100", 
"01000010110100001110010", "01000011001010110000000", "01000011100001010001110", "01000011110111110011100", 
"01000100001110010101100", "01000100100010110100000", "01000100111001010110000", "01000101001111110111110", 
"01000101100110011001100", "01000101111100111011010", "01000110010011011101000", "01000110101001111110110", 
"01000110111110011101100", "01000111010100111111010", "01000111101011100001010", "01001000000010000011000", 
"01001000011000100100110", "01001000101111000110100", "01001001000101101000010", "01001001011100001010000", 
"01001001110010101100000", "01001010000111001010110", "01001010011101101100100", "01001010110100001110010", 
"01001011001010110000000", "01001011100001010001110", "01001011110111110011100", "01001100001110010101100", 
"01001100100010110100000", "01001100111001010110000", "01001101001111110111110", "01001101100110011001100", 
"01001101111100111011010", "01001110010011011101000", "01001110101001111110110", "01001111000000100000110", 
"01001111010111000010100", "01001111101011100001010", "01010000000010000011000", "01010000011000100100110", 
"01010000101111000110100", "01010001000101101000010", "01010001011100001010000", "01010001110010101100000", 
"01010010001001001101110", "01010010011101101100100", "01010010110100001110010", "01010011001010110000000", 
"01010011100001010001110", "01010011110111110011100", "01010100001110010101100", "01010100100100110111010", 
"01010100111001010110000", "01010101001111110111110", "01010101100110011001100", "01010101111100111011010", 
"01010110010011011101000", "01010110101001111110110", "01010111000000100000110", "01010111010111000010100", 
"01010111101101100100010", "01011000000010000011000", "01011000011000100100110", "01011000101111000110100", 
"01011001000101101000010", "01011001011100001010000", "01011001110010101100000", "01011010001001001101110", 
"01011010011101101100100", "01011010110100001110010", "01011011001010110000000", "01011011100001010001110", 
"01011011110111110011100", "01011100001110010101100", "01011100100100110111010", "01011100111011011001000", 
"01011101010001111010110", "01011101100110011001100", "01011101111100111011010", "01011110010011011101000", 
"01011110101001111110110", "01011111000000100000110", "01011111010111000010100", "01011111101101100100010", 
"01100000000010000011000", "01100000011000100100110", "01100000101111000110100", "01100001000101101000010", 
"01100001011100001010000", "01100001110010101100000", "01100010001001001101110", "01100010011111101111100", 
"01100010110110010001010", "01100011001010110000000", "01100011100001010001110", "01100011110111110011100", 
"01100100001110010101100", "01100100100100110111010", "01100100111011011001000", "01100101010001111010110", 
"01100101101000011100100", "01100101111100111011010", "01100110010011011101000", "01100110101001111110110", 
"01100111000000100000110", "01100111010111000010100", "01100111101101100100010", "01101000000100000110000", 
"01101000011000100100110", "01101000101111000110100", "01101001000101101000010", "01101001011100001010000", 
"01101001110010101100000", "01101010001001001101110", "01101010011111101111100", "01101010110110010001010", 
"01101011001100110011000", "01101011100001010001110", "01101011110111110011100", "01101100001110010101100", 
"01101100100100110111010", "01101100111011011001000", "01101101010001111010110", "01101101101000011100100", 
"01101101111100111011010", "01101110010011011101000", "01101110101001111110110", "01101111000000100000110", 
"01101111010111000010100", "01101111101101100100010", "01110000000100000110000", "01110000011010100111110", 
"01110000110001001001100", "01110001000101101000010", "01110001011100001010000", "01110001110010101100000", 
"01110010001001001101110", "01110010011111101111100", "01110010110110010001010", "01110011001100110011000", 
"01110011100001010001110", "01110011110111110011100", "01110100001110010101100", "01110100100100110111010", 
"01110100111011011001000", "01110101010001111010110", "01110101101000011100100", "01110101111110111110010", 
"01110110010101100000010", "01110110101001111110110", "01110111000000100000110", "01110111010111000010100", 
"01110111101101100100010", "01111000000100000110000", "01111000011010100111110", "01111000110001001001100", 
"01111001000101101000010", "01111001011100001010000", "01111001110010101100000", "01111010001001001101110", 
"01111010011111101111100", "01111010110110010001010", "01111011001100110011000", "01111011100011010100110", 
"01111011110111110011100", "01111100001110010101100", "01111100100100110111010", "01111100111011011001000", 
"01111101010001111010110", "01111101101000011100100", "01111101111110111110010", "01111110010101100000010", 
"01111110101100000010000", "01111111000000100000110", "01111111010111000010100", "01111111101101100100010", 
"10000000000100000110000", "10000000011010100111110", "10000000110001001001100", "10000001000111101011100", 
"10000001011100001010000", "10000001110010101100000", "10000010001001001101110", "10000010011111101111100", 
"10000010110110010001010", "10000011001100110011000", "10000011100011010100110", "10000011111001110110110", 
"10000100001110010101100", "10000100100100110111010", "10000100111011011001000", "10000101010001111010110", 
"10000101101000011100100", "10000101111110111110010", "10000110010101100000010", "10000110101100000010000", 
"10000111000010100011110", "10000111010111000010100", "10000111101101100100010", "10001000000100000110000", 
"10001000011010100111110", "10001000110001001001100", "10001001000111101011100", "10001001011110001101010", 
"10001001110100101111000", "10001010001001001101110", "10001010011111101111100", "10001010110110010001010", 
"10001011001100110011000", "10001011100011010100110", "10001011111001110110110", "10001100010000011000100", 
"10001100100100110111010", "10001100111011011001000", "10001101010001111010110", "10001101101000011100100", 
"10001101111110111110010", "10001110010101100000010", "10001110101100000010000", "10001111000010100011110", 
"10001111010111000010100", "10001111101101100100010", "10010000000100000110000", "10010000011010100111110", 
"10010000110001001001100", "10010001000111101011100", "10010001011110001101010", "10010001110100101111000", 
"10010010001011010000110", "10010010011111101111100", "10010010110110010001010", "10010011001100110011000", 
"10010011100011010100110", "10010011111001110110110", "10010100010000011000100", "10010100100110111010010", 
"10010100111101011100000", "10010101010001111010110", "10010101101000011100100", "10010101111110111110010", 
"10010110010101100000010", "10010110101100000010000", "10010111000010100011110", "10010111011001000101100", 
"10010111101101100100010", "10011000000100000110000", "10011000011010100111110", "10011000110001001001100", 
"10011001000111101011100", "10011001011110001101010", "10011001110100101111000", "10011010001011010000110", 
"10011010100001110010100", "10011010110110010001010", "10011011001100110011000", "10011011100011010100110", 
"10011011111001110110110", "10011100010000011000100", "10011100100110111010010", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000"
);
type muon_muon_diff_phi_lut_ufixed_array is array (0 to 2**(MUON_PHI_HIGH-MUON_PHI_LOW+1)-1) of ufixed(2 downto -20);
constant MU_MU_DIFF_PHI_LUT_UFIXED : muon_muon_diff_phi_lut_ufixed_array := (
"00000000000000000000000", "00000000010110100001110", "00000000101101000011100", "00000001000011100101010", 
"00000001011010000111000", "00000001110000101000110", "00000010000101000111100", "00000010011011101001010", 
"00000010110010001011010", "00000011001000101101000", "00000011011111001110110", "00000011110101110000100", 
"00000100001100010010010", "00000100100010110100000", "00000100111001010110000", "00000101001111110111110", 
"00000101100110011001100", "00000101111010111000010", "00000110010001011010000", "00000110100111111011110", 
"00000110111110011101100", "00000111010100111111010", "00000111101011100001010", "00001000000010000011000", 
"00001000011000100100110", "00001000101111000110100", "00001001000101101000010", "00001001011100001010000", 
"00001001110000101000110", "00001010000111001010110", "00001010011101101100100", "00001010110100001110010", 
"00001011001010110000000", "00001011100001010001110", "00001011110111110011100", "00001100001110010101100", 
"00001100100100110111010", "00001100111011011001000", "00001101010001111010110", "00001101100110011001100", 
"00001101111100111011010", "00001110010011011101000", "00001110101001111110110", "00001111000000100000110", 
"00001111010111000010100", "00001111101101100100010", "00010000000100000110000", "00010000011010100111110", 
"00010000110001001001100", "00010001000111101011100", "00010001011100001010000", "00010001110010101100000", 
"00010010001001001101110", "00010010011111101111100", "00010010110110010001010", "00010011001100110011000", 
"00010011100011010100110", "00010011111001110110110", "00010100010000011000100", "00010100100110111010010", 
"00010100111011011001000", "00010101010001111010110", "00010101101000011100100", "00010101111110111110010", 
"00010110010101100000010", "00010110101100000010000", "00010111000010100011110", "00010111011001000101100", 
"00010111101111100111010", "00011000000110001001000", "00011000011100101011000", "00011000110001001001100", 
"00011001000111101011100", "00011001011110001101010", "00011001110100101111000", "00011010001011010000110", 
"00011010100001110010100", "00011010111000010100010", "00011011001110110110010", "00011011100101011000000", 
"00011011111011111001110", "00011100010010011011100", "00011100100110111010010", "00011100111101011100000", 
"00011101010011111101110", "00011101101010011111100", "00011110000001000001100", "00011110010111100011010", 
"00011110101110000101000", "00011111000100100110110", "00011111011011001000100", "00011111110001101010010", 
"00100000001000001100010", "00100000011100101011000", "00100000110011001100110", "00100001001001101110100", 
"00100001100000010000010", "00100001110110110010000", "00100010001101010011110", "00100010100011110101110", 
"00100010111010010111100", "00100011010000111001010", "00100011100111011011000", "00100011111101111100110", 
"00100100010010011011100", "00100100101000111101010", "00100100111111011111000", "00100101010110000001000", 
"00100101101100100010110", "00100110000011000100100", "00100110011001100110010", "00100110110000001000000", 
"00100111000110101001110", "00100111011101001011110", "00100111110011101101100", "00101000001000001100010", 
"00101000011110101110000", "00101000110101001111110", "00101001001011110001100", "00101001100010010011010", 
"00101001111000110101000", "00101010001111010111000", "00101010100101111000110", "00101010111100011010100", 
"00101011010010111100010", "00101011101001011110000", "00101011111101111100110", "00101100010100011110100", 
"00101100101011000000100", "00101101000001100010010", "00101101011000000100000", "00101101101110100101110", 
"00101110000101000111100", "00101110011011101001010", "00101110110010001011010", "00101111001000101101000", 
"00101111011111001110110", "00101111110011101101100", "00110000001010001111010", "00110000100000110001000", 
"00110000110111010010110", "00110001001101110100100", "00110001100100010110100", "00110001111010111000010", 
"00110010010001011010000", "00110010100111111011110", "00110010111110011101100", "00110011010100111111010", 
"00110011101001011110000", "00110011111111111111110", "00110100010110100001110", "00110100101101000011100", 
"00110101000011100101010", "00110101011010000111000", "00110101110000101000110", "00110110000111001010110", 
"00110110011101101100100", "00110110110100001110010", "00110111001010110000000", "00110111011111001110110", 
"00110111110101110000100", "00111000001100010010010", "00111000100010110100000", "00111000111001010110000", 
"00111001001111110111110", "00111001100110011001100", "00111001111100111011010", "00111010010011011101000", 
"00111010101001111110110", "00111011000000100000110", "00111011010100111111010", "00111011101011100001010", 
"00111100000010000011000", "00111100011000100100110", "00111100101111000110100", "00111101000101101000010", 
"00111101011100001010000", "00111101110010101100000", "00111110001001001101110", "00111110011111101111100", 
"00111110110100001110010", "00111111001010110000000", "00111111100001010001110", "00111111110111110011100", 
"01000000001110010101100", "01000000100100110111010", "01000000111011011001000", "01000001010001111010110", 
"01000001101000011100100", "01000001111110111110010", "01000010010101100000010", "01000010101001111110110", 
"01000011000000100000110", "01000011010111000010100", "01000011101101100100010", "01000100000100000110000", 
"01000100011010100111110", "01000100110001001001100", "01000101000111101011100", "01000101011110001101010", 
"01000101110100101111000", "01000110001011010000110", "01000110011111101111100", "01000110110110010001010", 
"01000111001100110011000", "01000111100011010100110", "01000111111001110110110", "01001000010000011000100", 
"01001000100110111010010", "01001000111101011100000", "01001001010011111101110", "01001001101010011111100", 
"01001010000001000001100", "01001010010101100000010", "01001010101100000010000", "01001011000010100011110", 
"01001011011001000101100", "01001011101111100111010", "01001100000110001001000", "01001100011100101011000", 
"01001100110011001100110", "01001101001001101110100", "01001101100000010000010", "01001101110110110010000", 
"01001110001011010000110", "01001110100001110010100", "01001110111000010100010", "01001111001110110110010", 
"01001111100101011000000", "01001111111011111001110", "01010000010010011011100", "01010000101000111101010", 
"01010000111111011111000", "01010001010110000001000", "01010001101100100010110", "01010010000001000001100", 
"01010010010111100011010", "01010010101110000101000", "01010011000100100110110", "01010011011011001000100", 
"01010011110001101010010", "01010100001000001100010", "01010100011110101110000", "01010100110101001111110", 
"01010101001011110001100", "01010101100010010011010", "01010101110110110010000", "01010110001101010011110", 
"01010110100011110101110", "01010110111010010111100", "01010111010000111001010", "01010111100111011011000", 
"01010111111101111100110", "01011000010100011110100", "01011000101011000000100", "01011001000001100010010", 
"01011001011000000100000", "01011001101100100010110", "01011010000011000100100", "01011010011001100110010", 
"01011010110000001000000", "01011011000110101001110", "01011011011101001011110", "01011011110011101101100", 
"01011100001010001111010", "01011100100000110001000", "01011100110111010010110", "01011101001101110100100", 
"01011101100010010011010", "01011101111000110101000", "01011110001111010111000", "01011110100101111000110", 
"01011110111100011010100", "01011111010010111100010", "01011111101001011110000", "01100000000000000000000", 
"01100000010110100001110", "01100000101101000011100", "01100001000011100101010", "01100001011000000100000", 
"01100001101110100101110", "01100010000101000111100", "01100010011011101001010", "01100010110010001011010", 
"01100011001000101101000", "01100011011111001110110", "01100011110101110000100", "01100100001100010010010", 
"01100100100010110100000", "01100100111001010110000", "01100101001101110100100", "01100101100100010110100", 
"01100101111010111000010", "01100110010001011010000", "01100110100111111011110", "01100110111110011101100", 
"01100111010100111111010", "01100111101011100001010", "01101000000010000011000", "01101000011000100100110", 
"01101000101101000011100", "01101001000011100101010", "01101001011010000111000", "01101001110000101000110", 
"01101010000111001010110", "01101010011101101100100", "01101010110100001110010", "01101011001010110000000", 
"01101011100001010001110", "01101011110111110011100", "01101100001110010101100", "01101100100010110100000", 
"01101100111001010110000", "01101101001111110111110", "01101101100110011001100", "01101101111100111011010", 
"01101110010011011101000", "01101110101001111110110", "01101111000000100000110", "01101111010111000010100", 
"01101111101101100100010", "01110000000100000110000", "01110000011000100100110", "01110000101111000110100", 
"01110001000101101000010", "01110001011100001010000", "01110001110010101100000", "01110010001001001101110", 
"01110010011111101111100", "01110010110110010001010", "01110011001100110011000", "01110011100011010100110", 
"01110011111001110110110", "01110100001110010101100", "01110100100100110111010", "01110100111011011001000", 
"01110101010001111010110", "01110101101000011100100", "01110101111110111110010", "01110110010101100000010", 
"01110110101100000010000", "01110111000010100011110", "01110111011001000101100", "01110111101111100111010", 
"01111000000100000110000", "01111000011010100111110", "01111000110001001001100", "01111001000111101011100", 
"01111001011110001101010", "01111001110100101111000", "01111010001011010000110", "01111010100001110010100", 
"01111010111000010100010", "01111011001110110110010", "01111011100101011000000", "01111011111001110110110", 
"01111100010000011000100", "01111100100110111010010", "01111100111101011100000", "01111101010011111101110", 
"01111101101010011111100", "01111110000001000001100", "01111110010111100011010", "01111110101110000101000", 
"01111111000100100110110", "01111111011011001000100", "01111111101111100111010", "10000000000110001001000", 
"10000000011100101011000", "10000000110011001100110", "10000001001001101110100", "10000001100000010000010", 
"10000001110110110010000", "10000010001101010011110", "10000010100011110101110", "10000010111010010111100", 
"10000011010000111001010", "10000011100101011000000", "10000011111011111001110", "10000100010010011011100", 
"10000100101000111101010", "10000100111111011111000", "10000101010110000001000", "10000101101100100010110", 
"10000110000011000100100", "10000110011001100110010", "10000110110000001000000", "10000111000110101001110", 
"10000111011011001000100", "10000111110001101010010", "10001000001000001100010", "10001000011110101110000", 
"10001000110101001111110", "10001001001011110001100", "10001001100010010011010", "10001001111000110101000", 
"10001010001111010111000", "10001010100101111000110", "10001010111100011010100", "10001011010000111001010", 
"10001011100111011011000", "10001011111101111100110", "10001100010100011110100", "10001100101011000000100", 
"10001101000001100010010", "10001101011000000100000", "10001101101110100101110", "10001110000101000111100", 
"10001110011011101001010", "10001110110000001000000", "10001111000110101001110", "10001111011101001011110", 
"10001111110011101101100", "10010000001010001111010", "10010000100000110001000", "10010000110111010010110", 
"10010001001101110100100", "10010001100100010110100", "10010001111010111000010", "10010010010001011010000", 
"10010010100101111000110", "10010010111100011010100", "10010011010010111100010", "10010011101001011110000", 
"10010011111111111111110", "10010100010110100001110", "10010100101101000011100", "10010101000011100101010", 
"10010101011010000111000", "10010101110000101000110", "10010110000111001010110", "10010110011011101001010", 
"10010110110010001011010", "10010111001000101101000", "10010111011111001110110", "10010111110101110000100", 
"10011000001100010010010", "10011000100010110100000", "10011000111001010110000", "10011001001111110111110", 
"10011001100110011001100", "10011001111100111011010", "10011010010001011010000", "10011010100111111011110", 
"10011010111110011101100", "10011011010100111111010", "10011011101011100001010", "10011100000010000011000", 
"10011100011000100100110", "10011100101111000110100", "10011101000101101000010", "10011101011100001010000", 
"10011101110010101100000", "10011110000111001010110", "10011110011101101100100", "10011110110100001110010", 
"10011111001010110000000", "10011111100001010001110", "10011111110111110011100", "10100000001110010101100", 
"10100000100100110111010", "10100000111011011001000", "10100001010001111010110", "10100001101000011100100", 
"10100001111100111011010", "10100010010011011101000", "10100010101001111110110", "10100011000000100000110", 
"10100011010111000010100", "10100011101101100100010", "10100100000100000110000", "10100100011010100111110", 
"10100100110001001001100", "10100101000111101011100", "10100101011110001101010", "10100101110010101100000", 
"10100110001001001101110", "10100110011111101111100", "10100110110110010001010", "10100111001100110011000", 
"10100111100011010100110", "10100111111001110110110", "10101000010000011000100", "10101000100110111010010", 
"10101000111101011100000", "10101001010011111101110", "10101001101000011100100", "10101001111110111110010", 
"10101010010101100000010", "10101010101100000010000", "10101011000010100011110", "10101011011001000101100", 
"10101011101111100111010", "10101100000110001001000", "10101100011100101011000", "10101100110011001100110", 
"10101101001001101110100", "10101101011110001101010", "10101101110100101111000", "10101110001011010000110", 
"10101110100001110010100", "10101110111000010100010", "10101111001110110110010", "10101111100101011000000", 
"10101111111011111001110", "10110000010010011011100", "10110000101000111101010", "10110000111111011111000", 
"10110001010011111101110", "10110001101010011111100", "10110010000001000001100", "10110010010111100011010", 
"10110010101110000101000", "10110011000100100110110", "10110011011011001000100", "10110011110001101010010", 
"10110100001000001100010", "10110100011110101110000", "10110100110101001111110", "10110101001001101110100", 
"10110101100000010000010", "10110101110110110010000", "10110110001101010011110", "10110110100011110101110", 
"10110110111010010111100", "10110111010000111001010", "10110111100111011011000", "10110111111101111100110", 
"10111000010100011110100", "10111000101000111101010", "10111000111111011111000", "10111001010110000001000", 
"10111001101100100010110", "10111010000011000100100", "10111010011001100110010", "10111010110000001000000", 
"10111011000110101001110", "10111011011101001011110", "10111011110011101101100", "10111100001010001111010", 
"10111100011110101110000", "10111100110101001111110", "10111101001011110001100", "10111101100010010011010", 
"10111101111000110101000", "10111110001111010111000", "10111110100101111000110", "10111110111100011010100", 
"10111111010010111100010", "10111111101001011110000", "11000000000000000000000", "11000000010100011110100", 
"11000000101011000000100", "11000001000001100010010", "11000001011000000100000", "11000001101110100101110", 
"11000010000101000111100", "11000010011011101001010", "11000010110010001011010", "11000011001000101101000", 
"11000011011111001110110", "11000011110101110000100", "11000100001010001111010", "11000100100000110001000", 
"11000100110111010010110", "11000101001101110100100", "11000101100100010110100", "11000101111010111000010", 
"11000110010001011010000", "11000110100111111011110", "11000110111110011101100", "11000111010100111111010", 
"11000111101011100001010", "11000111111111111111110", "11001000010110100001110", "11001000101101000011100", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000", 
"00000000000000000000000", "00000000000000000000000", "00000000000000000000000", "00000000000000000000000"
);
type muon_muon_cosh_deta_lut_ufixed_array is array (0 to 2**(MUON_ETA_HIGH-MUON_ETA_LOW+1)-1) of ufixed(6 downto -20);
constant MU_MU_COSH_DETA_LUT_UFIXED : muon_muon_cosh_deta_lut_ufixed_array := (
"000000100000000000000000000", "000000100000000000001101000", "000000100000000000011010000", "000000100000000001000001100", 
"000000100000000001110101110", "000000100000000011000100100", "000000100000000100010011010", "000000100000000101111100000", 
"000000100000000111110010000", "000000100000001001110101000", "000000100000001100000101010", "000000100000001110101111100", 
"000000100000010001011010000", "000000100000010100011110100", "000000100000010111110000010", "000000100000011011001111010", 
"000000100000011111001000010", "000000100000100011000001010", "000000100000100111010100100", "000000100000101011110100110", 
"000000100000110000100010010", "000000100000110101101010000", "000000100000111010111110110", "000000100001000000010011100", 
"000000100001000110001111110", "000000100001001100001011110", "000000100001010010010101000", "000000100001011000111000100", 
"000000100001011111101001000", "000000100001100110100110100", "000000100001101101111110100", "000000100001110101100011100", 
"000000100001111101010101100", "000000100010000101010100110", "000000100010001101100001000", "000000100010010110000111100", 
"000000100010011110111011000", "000000100010101000001001000", "000000100010110001010110110", "000000100010111010111110110", 
"000000100011000100110100000", "000000100011001111000011010", "000000100011011001010010100", "000000100011100011111100010", 
"000000100011101111000000000", "000000100011111010010000110", "000000100100000101101111000", "000000100100010001011010000", 
"000000100100011101011111010", "000000100100101001110001110", "000000100100110110010001010", "000000100101000011001011000", 
"000000100101010000010010000", "000000100101011101110011000", "000000100101101011010100000", "000000100101111001011100100", 
"000000100110000111100100110", "000000100110010110010100100", "000000100110100101000100010", "000000100110110100001110010", 
"000000100111000011100101010", "000000100111010011010110100", "000000100111100011010100110", "000000100111110011101101100", 
"000000101000000100010011010", "000000101000010101010011000", "000000101000100110100000000", "000000101000111000000111010", 
"000000101001001001111011100", "000000101001011100001010000", "000000101001101110100101110", "000000101010000001011011110", 
"000000101010010100011110100", "000000101010100111111011110", "000000101010111011110011010", "000000101011001111110111110", 
"000000101011100100001001010", "000000101011111001000010010", "000000101100001110001000010", "000000101100100011011011100", 
"000000101100111001001000110", "000000101101001111010000010", "000000101101100101110010010", "000000101101111100100001000", 
"000000101110010011101010010", "000000101110101011000000100", "000000101111000010111110000", "000000101111011011001000100", 
"000000101111110011101101100", "000000110000001100011111100", "000000110000100101111000110", "000000110000111111011111000", 
"000000110001011001011111110", "000000110001110011101101100", "000000110010001110100010100", "000000110010101001110001110", 
"000000110011000101001110000", "000000110011100001000100110", "000000110011111101010101100", "000000110100011010001101100", 
"000000110100110111010010110", "000000110101010100110010010", "000000110101110010011110110", "000000110110010000110010110", 
"000000110110101111100000110", "000000110111001110101001000", "000000110111101110001011100", "000000111000001110001000010", 
"000000111000101110011111010", "000000111001001111011101100", "000000111001110000101000110", "000000111010010010011011100", 
"000000111010110100011011010", "000000111011010111000010100", "000000111011111010000011110", "000000111100011101011111010", 
"000000111101000001100010010", "000000111101100101110010010", "000000111110001010101001100", "000000111110110000001000000", 
"000000111111010101110011110", "000000111111111100000110110", "000001000000100011000001010", "000001000001001010001000110", 
"000001000001110001110111100", "000001000010011010001101100", "000001000011000010111110000", "000001000011101100001000100", 
"000001000100010101111010010", "000001000101000000010011100", "000001000101101011000111000", "000001000110010110010100100", 
"000001000111000010010110100", "000001000111101110110010110", "000001001000011011101001010", "000001001001001001000111010", 
"000001001001110111001100010", "000001001010100101111000110", "000001001011010100111111010", "000001001100000100101101010", 
"000001001100110101000010110", "000001001101100101111111010", "000001001110010111100011010", "000001001111001001100001010", 
"000001001111111100010100000", "000001010000101111100000110", "000001010001100011100010000", "000001010010010111111101100", 
"000001010011001101000000010", "000001010100000010110111100", "000001010100111001010110000", "000001010101110000011011110", 
"000001010110100111111011110", "000001010111100000011101010", "000001011000011001011001010", "000001011001010011001001100", 
"000001011010001101100001000", "000001011011001000011111110", "000001011100000100010011010", "000001011101000000101101110", 
"000001011101111101101111110", "000001011110111011100110000", "000001011111111010010000110", "000001100000111001100011000", 
"000001100001111001011100100", "000001100010111010010111100", "000001100011111011111001110", "000001100100111110000011010", 
"000001100110000001001110100", "000001100111000101000001000", "000001101000001001101000000", "000001101001001110110110010", 
"000001101010010101000110000", "000001101011011100001010000", "000001101100100011110101110", "000001101101101100100010110", 
"000001101110110101110111000", "000001110000000000001101000", "000001110001001011010111010", "000001110010010111010110000", 
"000001110011100100001001010", "000001110100110001111110000", "000001110110000000011010000", "000001110111010000000100110", 
"000001111000100000010110110", "000001111001110001101010010", "000001111011000011111111100", "000001111100010111001001000", 
"000001111101101011010100000", "000001111111000000010011100", "000010000000010110010100100", "000010000001101101010111000", 
"000010000011000101001110000", "000010000100011110010011110", "000010000101111000001101110", "000010000111010011010110100", 
"000010001000101111010011110", "000010001010001100010010010", "000010001011101010011111100", "000010001101001001100001010", 
"000010001110101001110001110", "000010010000001011000011110", "000010010001101101010111000", "000010010011010000111001010", 
"000010010100110101101010000", "000010010110011011001111010", "000010011000000010010000000", "000010011001101010000101100", 
"000010011011010011010110100", "000010011100111101101001010", "000010011110101001010111100", "000010100000010110000111100", 
"000010100010000100000110000", "000010100011110011000110000", "000010100101100011100010000", "000010100111010101001100100", 
"000010101001001000010010110", "000010101010111100011010100", "000010101100110001111110000", "000010101110101000110000010", 
"000010110000100000111110010", "000010110010011010011010110", "000010110100010101010011000", "000010110110010001100111000", 
"000010111000001111001001110", "000010111010001110001000010", "000010111100001110100010100", "000010111110010000011000100", 
"000011000000010011011101000", "000011000010011000001010100", "000011000100011110100000110", "000011000110100110000101110", 
"000011001000101111010011110", "000011001010111001111101010", "000011001101000110001111110", "000011001111010011111101110", 
"000011010001100011010100110", "000011010011110100010100110", "000011010110000110110000100", "000011011000011011000010000", 
"000011011010110000101111100", "000011011101001000000101100", "000011011111100001010001110", "000011100001111100000110110", 
"000011100100011000100100110", "000011100110110110111000100", "000011101001010110110101010", "000011101011111000101000000", 
"000011101110011100010000110", "000011110001000001100010010", "000011110011101000110110110", "000011110110010001110100010", 
"000011111000111100100111100", "000011111011101001011110000", "000011111110011000001010100", "000100000001001000101101000", 
"000100000011111011010010100", "000100000110101111111011000", "000100001001100110011001100", "000100001100011110111011000", 
"000100001111011001011111110", "000100010010010101111010010", "000100010101010100110010010", "000100011000010101100000010", 
"000100011011011000011110010", "000100011110011101011111010", "000100100001100100100011100", "000100100100101110000101000", 
"000100100111111001101001100", "000100101011000111011110010", "000100101110010111110000010", "000100110001101010000101100", 
"000100110100111110110111110", "000100111000010101111010010", "000100111011101111011010010", "000100111111001011001010010", 
"000101000010101001010111100", "000101000110001010000010010", "000101001001101101001010000", "000101001101010010111100010", 
"000101010000111010111110110", "000101010100100101101011100", "000101011000010011000010110", "000101011100000010110111100", 
"000101011111110101100011100", "000101100011101010101100110", "000101100111100010100000100", "000101101011011101001011110", 
"000101101111011010100001010", "000101110011011010101110010", "000101110111011101100101110", "000101111011100011010100110", 
"000101111111101100001000100", "000110000011110111100110100", "000110001000000110001001000", "000110001100010111110000010", 
"000110010000101100000010000", "000110010101000011100101010", "000110011001011110001101010", "000110011101111011111001110", 
"000110100010011100101011000", "000110100111000000101101110", "000110101011100111110101010", "000110110000010010001110100", 
"000110110100111111111001010", "000110111001110001000011000", "000110111110100101010001100", "000111000011011100111110100", 
"000111001000011000001010100", "000111001101010110110101010", "000111010010011000110001110", "000111010111011110011010010", 
"000111011100100111100001100", "000111100001110100010100110", "000111100111000100110100000", "000111101100011000111111000", 
"000111110001110000110110000", "000111110111001100011000110", "000111111100101011110100110", "001000000010001111001001110", 
"001000000111110110010111110", "001000001101100001011111000", "001000010011010000011111000", "001000011001000011100101010", 
"001000011110111010110001110", "001000100100110110000100010", "001000101010110101011100110", "001000110000111001001000110", 
"001000110111000000111010110", "001000111101001101001101010", "001001000011011101100101110", "001001001001110010011110110", 
"001001010000001011111000000", "001001010110101001100100110", "001001011101001011111110110", "001001100011110010111001000", 
"001001101010011110100000110", "001001110001001110101001000", "001001111000000011101011110", "001001111110111101011100000", 
"001010000101111011111001110", "001010001100111111011111000", "001010010100000111111111000", "001010011011010101011001100", 
"001010100010100111101110110", "001010101001111111011000100", "001010110001011100001010000", "001010111000111110000011010", 
"001011000000100101010001100", "001011001000010001110100010", "001011010000000011101011110", "001011010111111011000101010", 
"001011011111111000000000110", "001011100111111010011110000", "001011110000000010101010010", "001011111000010000011000100", 
"001100000000100100000010110", "001100001000111101011100000", "001100010001011100100100010", "001100011010000001110101110", 
"001100100010101101000011100", "001100101011011110011010010", "001100110100010101101101010", "001100111101010011010110100", 
"001101000110010111010110000", "001101001111100001101100000", "001101011000110010001011010", "001101100010001001011010110", 
"001101101011100111001110000", "001101110101001011100100100", "001101111110110110011110100", "001110001000101000010110000", 
"001110010010100000111110010", "001110011100100000100100000", "001110100110100111000111010", "001110110000110100110101100", 
"001110111011001001101110100", "001111000101100101110010010", "001111010000001001000000100", "001111011010110011110100000", 
"001111100101100101111111010", "001111110000011111101111100", "001111111011100001000100110", "010000000110101010001100000", 
"010000010001111011000101010", "010000011101010011111101110", "010000101000110100101000100", "010000110100011101011111010", 
"010001000000001110100010100", "010001001100000111110010000", "010001011000001001001101110", "010001100100010011010000000", 
"010001110000100101101011100", "010001111101000000101101110", "010010001001100100100011100", "010010010110010000111111110", 
"010010100011000110011100110", "010010110000000100111010100", "010010111101001100011000110", "010011001010011101000101000", 
"010011010111110111001100010", "010011100101011010100001010", "010011110011000111011110010", "010100000000111101110110010", 
"010100001110111110000011010", "010100011101000111111000100", "010100101011011011110000000", "010100111001111001101001100", 
"010101001000100001100101100", "010101010111010011110000110", "010101100110010000011000100", "010101110101010111011100110", 
"010110000100101001001010100", "010110010100000101010100110", "010110100011101100100010110", "010110110011011110100111100", 
"010111000011011011110000000", "010111010011100011111100010", "010111100011110111011001010", "010111110100010110100001110", 
"011000000101000000111010110", "011000010101110111001100010", "011000100110111001001000110", "011000111000000110111101100", 
"011001001001100000110111100", "011001011011000111000100000", "011001101100111001010110000", "011001111110111000010100010", 
"011010010001000011110010010", "011010100011011011111101000", "011010110110000001000001100", "011011001000110010111111100", 
"011011011011110010010001110", "011011101110111110110111110", "011100000010011000110001110", "011100010110000000001101000", 
"011100101001110101100011100", "011100111101111000101000000", "011101010010001001110101000", "011101100110101001001010100", 
"011101111011010110110101010", "011110010000010010110101110", "011110100101011101110011000", "011110111010110111100000000", 
"011111010000011111111100100", "011111100110010111110000010", "011111111100011110111011000", "100000010010110101011100110", 
"100000101001011011100010110", "100001000000010001100111000", "100001010111010111101001110", "000000000000000000000000000", 
"000000000000000000000000000", "000000000000000000000000000", "000000000000000000000000000", "000000000000000000000000000", 
"000000000000000000000000000", "000000000000000000000000000", "000000000000000000000000000", "000000000000000000000000000", 
"000000000000000000000000000", "000000000000000000000000000", "000000000000000000000000000", "000000000000000000000000000", 
"000000000000000000000000000", "000000000000000000000000000", "000000000000000000000000000", "000000000000000000000000000", 
"000000000000000000000000000", "000000000000000000000000000", "000000000000000000000000000", "000000000000000000000000000", 
"000000000000000000000000000", "000000000000000000000000000", "000000000000000000000000000", "000000000000000000000000000", 
"000000000000000000000000000", "000000000000000000000000000", "000000000000000000000000000", "000000000000000000000000000", 
"000000000000000000000000000", "000000000000000000000000000", "000000000000000000000000000", "000000000000000000000000000", 
"000000000000000000000000000", "000000000000000000000000000", "000000000000000000000000000", "000000000000000000000000000", 
"000000000000000000000000000", "000000000000000000000000000", "000000000000000000000000000", "000000000000000000000000000", 
"000000000000000000000000000", "000000000000000000000000000", "000000000000000000000000000", "000000000000000000000000000", 
"000000000000000000000000000", "000000000000000000000000000", "000000000000000000000000000", "000000000000000000000000000", 
"000000000000000000000000000", "000000000000000000000000000", "000000000000000000000000000", "000000000000000000000000000", 
"000000000000000000000000000", "000000000000000000000000000", "000000000000000000000000000", "000000000000000000000000000", 
"000000000000000000000000000", "000000000000000000000000000", "000000000000000000000000000", "000000000000000000000000000"
);
type muon_muon_cos_dphi_lut_ufixed_array is array (0 to 2**(MUON_PHI_HIGH-MUON_PHI_LOW+1)-1) of ufixed(0 downto -20);
constant MU_MU_COS_DPHI_LUT_UFIXED : muon_muon_cos_dphi_lut_ufixed_array := (
"100000000000000000000", "011111111111110010110", "011111111111100101110", "011111111110111110010", 
"011111111101111100110", "011111111100111011010", "011111111011101100100", "011111111010000011110", 
"011111111000001101110", "011111110110001010110", "011111110011111010100", "011111110001010000010", 
"011111101110011000110", "011111101011100001010", "011111101000001111100", "011111100100100011100", 
"011111100000110111100", "011111011100111110100", "011111011000101011010", "011111010100001011000", 
"011111001111011101100", "011111001010100011000", "011111000101001110000", "011110111111111001010", 
"011110111010001010010", "011110110100001110010", "011110101110000101000", "011110100111101110110", 
"011110100001001011010", "011110011010011010110", "011110010011010000000", "011110001100000101010", 
"011110000100100000010", "011101111100101110010", "011101110100101111000", "011101101100100010110", 
"011101100100001001010", "011101011011100010110", "011101010010100010000", "011101001001100001010", 
"011101000000000110100", "011100110110011110100", "011100101100110110010", "011100100010110100000", 
"011100011000100100110", "011100001110001000010", "011100000011011110110", "011011111000101000000", 
"011011101101100100010", "011011100010010011010", "011011010110110101010", "011011001011001010010", 
"011010111111010010000", "011010110011001100110", "011010100110111010010", "011010011010011010110", 
"011010001101101110000", "011010000000100111010", "011001110011100000010", "011001100110001100010", 
"011001011000111000100", "011001001011001010010", "011000111101001111000", "011000101111000110100", 
"011000100000110001000", "011000010010011011100", "011000000011101011110", "010111110100111100000", 
"010111100101111111010", "010111010110110101010", "010111000111011110010", "010110110111111010010", 
"010110101000001001000", "010110011000010111110", "010110001000001100010", "010101111000000000110", 
"010101100111101000000", "010101010111000010100", "010101000110001111110", "010100110101011100110", 
"010100100100011101000", "010100010011010000000", "010100000001110101110", "010011110000011011110", 
"010011011110110100100", "010011001101000000010", "010010111010111110110", "010010101000111101010", 
"010010010110101110110", "010010000100010011010", "010001110001110111100", "010001011111001110110", 
"010001001100011000110", "010000111001100011000", "010000100110100000000", "010000010011010000000", 
"001111111111111111110", "001111101100100010110", "001111011001000101100", "001111000101011011010", 
"001110110001100011110", "001110011101101100100", "001110001001110101000", "001101110101110000100", 
"001101100001011111000", "001101001101001101010", "001100111000101110100", "001100100100001111110", 
"001100001111110001010", "001011111011000101010", "001011100110001100010", "001011010001100000100", 
"001010111100011010100", "001010100111010100100", "001010010010001110100", "001001111101001000010", 
"001001100111110101010", "001001010010100010000", "001000111101000001110", "001000100111100001100", 
"001000010010000001010", "000111111100100001000", "000111100110110011110", "000111010001000110010", 
"000110111011001011110", "000110100101011110100", "000110001111100100000", "000101111001101001100", 
"000101100011100010000", "000101001101100111100", "000100110111100000000", "000100100001011000010", 
"000100001011010000110", "000011110101001001010", "000011011111000001100", "000011001000101101000", 
"000010110010100101010", "000010011100010000110", "000010000101111100000", "000001101111100111010", 
"000001011001010010100", "000001000010111110000", "000000101100101001010", "000000010110010100100", 
"000000000000000000000", "000000010110010100100", "000000101100101001010", "000001000010111110000", 
"000001011001010010100", "000001101111100111010", "000010000101111100000", "000010011100010000110", 
"000010110010100101010", "000011001000101101000", "000011011111000001100", "000011110101001001010", 
"000100001011010000110", "000100100001011000010", "000100110111100000000", "000101001101100111100", 
"000101100011100010000", "000101111001101001100", "000110001111100100000", "000110100101011110100", 
"000110111011001011110", "000111010001000110010", "000111100110110011110", "000111111100100001000", 
"001000010010000001010", "001000100111100001100", "001000111101000001110", "001001010010100010000", 
"001001100111110101010", "001001111101001000010", "001010010010001110100", "001010100111010100100", 
"001010111100011010100", "001011010001100000100", "001011100110001100010", "001011111011000101010", 
"001100001111110001010", "001100100100001111110", "001100111000101110100", "001101001101001101010", 
"001101100001011111000", "001101110101110000100", "001110001001110101000", "001110011101101100100", 
"001110110001100011110", "001111000101011011010", "001111011001000101100", "001111101100100010110", 
"001111111111111111110", "010000010011010000000", "010000100110100000000", "010000111001100011000", 
"010001001100011000110", "010001011111001110110", "010001110001110111100", "010010000100010011010", 
"010010010110101110110", "010010101000111101010", "010010111010111110110", "010011001101000000010", 
"010011011110110100100", "010011110000011011110", "010100000001110101110", "010100010011010000000", 
"010100100100011101000", "010100110101011100110", "010101000110001111110", "010101010111000010100", 
"010101100111101000000", "010101111000000000110", "010110001000001100010", "010110011000010111110", 
"010110101000001001000", "010110110111111010010", "010111000111011110010", "010111010110110101010", 
"010111100101111111010", "010111110100111100000", "011000000011101011110", "011000010010011011100", 
"011000100000110001000", "011000101111000110100", "011000111101001111000", "011001001011001010010", 
"011001011000111000100", "011001100110001100010", "011001110011100000010", "011010000000100111010", 
"011010001101101110000", "011010011010011010110", "011010100110111010010", "011010110011001100110", 
"011010111111010010000", "011011001011001010010", "011011010110110101010", "011011100010010011010", 
"011011101101100100010", "011011111000101000000", "011100000011011110110", "011100001110001000010", 
"011100011000100100110", "011100100010110100000", "011100101100110110010", "011100110110011110100", 
"011101000000000110100", "011101001001100001010", "011101010010100010000", "011101011011100010110", 
"011101100100001001010", "011101101100100010110", "011101110100101111000", "011101111100101110010", 
"011110000100100000010", "011110001100000101010", "011110010011010000000", "011110011010011010110", 
"011110100001001011010", "011110100111101110110", "011110101110000101000", "011110110100001110010", 
"011110111010001010010", "011110111111111001010", "011111000101001110000", "011111001010100011000", 
"011111001111011101100", "011111010100001011000", "011111011000101011010", "011111011100111110100", 
"011111100000110111100", "011111100100100011100", "011111101000001111100", "011111101011100001010", 
"011111101110011000110", "011111110001010000010", "011111110011111010100", "011111110110001010110", 
"011111111000001101110", "011111111010000011110", "011111111011101100100", "011111111100111011010", 
"011111111101111100110", "011111111110111110010", "011111111111100101110", "011111111111110010110", 
"100000000000000000000", "011111111111110010110", "011111111111100101110", "011111111110111110010", 
"011111111101111100110", "011111111100111011010", "011111111011101100100", "011111111010000011110", 
"011111111000001101110", "011111110110001010110", "011111110011111010100", "011111110001010000010", 
"011111101110011000110", "011111101011100001010", "011111101000001111100", "011111100100100011100", 
"011111100000110111100", "011111011100111110100", "011111011000101011010", "011111010100001011000", 
"011111001111011101100", "011111001010100011000", "011111000101001110000", "011110111111111001010", 
"011110111010001010010", "011110110100001110010", "011110101110000101000", "011110100111101110110", 
"011110100001001011010", "011110011010011010110", "011110010011010000000", "011110001100000101010", 
"011110000100100000010", "011101111100101110010", "011101110100101111000", "011101101100100010110", 
"011101100100001001010", "011101011011100010110", "011101010010100010000", "011101001001100001010", 
"011101000000000110100", "011100110110011110100", "011100101100110110010", "011100100010110100000", 
"011100011000100100110", "011100001110001000010", "011100000011011110110", "011011111000101000000", 
"011011101101100100010", "011011100010010011010", "011011010110110101010", "011011001011001010010", 
"011010111111010010000", "011010110011001100110", "011010100110111010010", "011010011010011010110", 
"011010001101101110000", "011010000000100111010", "011001110011100000010", "011001100110001100010", 
"011001011000111000100", "011001001011001010010", "011000111101001111000", "011000101111000110100", 
"011000100000110001000", "011000010010011011100", "011000000011101011110", "010111110100111100000", 
"010111100101111111010", "010111010110110101010", "010111000111011110010", "010110110111111010010", 
"010110101000001001000", "010110011000010111110", "010110001000001100010", "010101111000000000110", 
"010101100111101000000", "010101010111000010100", "010101000110001111110", "010100110101011100110", 
"010100100100011101000", "010100010011010000000", "010100000001110101110", "010011110000011011110", 
"010011011110110100100", "010011001101000000010", "010010111010111110110", "010010101000111101010", 
"010010010110101110110", "010010000100010011010", "010001110001110111100", "010001011111001110110", 
"010001001100011000110", "010000111001100011000", "010000100110100000000", "010000010011010000000", 
"001111111111111111110", "001111101100100010110", "001111011001000101100", "001111000101011011010", 
"001110110001100011110", "001110011101101100100", "001110001001110101000", "001101110101110000100", 
"001101100001011111000", "001101001101001101010", "001100111000101110100", "001100100100001111110", 
"001100001111110001010", "001011111011000101010", "001011100110001100010", "001011010001100000100", 
"001010111100011010100", "001010100111010100100", "001010010010001110100", "001001111101001000010", 
"001001100111110101010", "001001010010100010000", "001000111101000001110", "001000100111100001100", 
"001000010010000001010", "000111111100100001000", "000111100110110011110", "000111010001000110010", 
"000110111011001011110", "000110100101011110100", "000110001111100100000", "000101111001101001100", 
"000101100011100010000", "000101001101100111100", "000100110111100000000", "000100100001011000010", 
"000100001011010000110", "000011110101001001010", "000011011111000001100", "000011001000101101000", 
"000010110010100101010", "000010011100010000110", "000010000101111100000", "000001101111100111010", 
"000001011001010010100", "000001000010111110000", "000000101100101001010", "000000010110010100100", 
"000000000000000000000", "000000010110010100100", "000000101100101001010", "000001000010111110000", 
"000001011001010010100", "000001101111100111010", "000010000101111100000", "000010011100010000110", 
"000010110010100101010", "000011001000101101000", "000011011111000001100", "000011110101001001010", 
"000100001011010000110", "000100100001011000010", "000100110111100000000", "000101001101100111100", 
"000101100011100010000", "000101111001101001100", "000110001111100100000", "000110100101011110100", 
"000110111011001011110", "000111010001000110010", "000111100110110011110", "000111111100100001000", 
"001000010010000001010", "001000100111100001100", "001000111101000001110", "001001010010100010000", 
"001001100111110101010", "001001111101001000010", "001010010010001110100", "001010100111010100100", 
"001010111100011010100", "001011010001100000100", "001011100110001100010", "001011111011000101010", 
"001100001111110001010", "001100100100001111110", "001100111000101110100", "001101001101001101010", 
"001101100001011111000", "001101110101110000100", "001110001001110101000", "001110011101101100100", 
"001110110001100011110", "001111000101011011010", "001111011001000101100", "001111101100100010110", 
"001111111111111111110", "010000010011010000000", "010000100110100000000", "010000111001100011000", 
"010001001100011000110", "010001011111001110110", "010001110001110111100", "010010000100010011010", 
"010010010110101110110", "010010101000111101010", "010010111010111110110", "010011001101000000010", 
"010011011110110100100", "010011110000011011110", "010100000001110101110", "010100010011010000000", 
"010100100100011101000", "010100110101011100110", "010101000110001111110", "010101010111000010100", 
"010101100111101000000", "010101111000000000110", "010110001000001100010", "010110011000010111110", 
"010110101000001001000", "010110110111111010010", "010111000111011110010", "010111010110110101010", 
"010111100101111111010", "010111110100111100000", "011000000011101011110", "011000010010011011100", 
"011000100000110001000", "011000101111000110100", "011000111101001111000", "011001001011001010010", 
"011001011000111000100", "011001100110001100010", "011001110011100000010", "011010000000100111010", 
"011010001101101110000", "011010011010011010110", "011010100110111010010", "011010110011001100110", 
"011010111111010010000", "011011001011001010010", "011011010110110101010", "011011100010010011010", 
"011011101101100100010", "011011111000101000000", "011100000011011110110", "011100001110001000010", 
"011100011000100100110", "011100100010110100000", "011100101100110110010", "011100110110011110100", 
"011101000000000110100", "011101001001100001010", "011101010010100010000", "011101011011100010110", 
"011101100100001001010", "011101101100100010110", "011101110100101111000", "011101111100101110010", 
"011110000100100000010", "011110001100000101010", "011110010011010000000", "011110011010011010110", 
"011110100001001011010", "011110100111101110110", "011110101110000101000", "011110110100001110010", 
"011110111010001010010", "011110111111111001010", "011111000101001110000", "011111001010100011000", 
"011111001111011101100", "011111010100001011000", "011111011000101011010", "011111011100111110100", 
"011111100000110111100", "011111100100100011100", "011111101000001111100", "011111101011100001010", 
"011111101110011000110", "011111110001010000010", "011111110011111010100", "011111110110001010110", 
"011111111000001101110", "011111111010000011110", "011111111011101100100", "011111111100111011010", 
"011111111101111100110", "011111111110111110010", "011111111111100101110", "011111111111110010110", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000", 
"000000000000000000000", "000000000000000000000", "000000000000000000000", "000000000000000000000"
);
type muon_muon_cos_dphi_sign_lut_array is array (0 to 2**(MUON_PHI_HIGH-MUON_PHI_LOW+1)-1) of boolean;
constant MU_MU_COS_DPHI_SIGN_LUT : muon_muon_cos_dphi_sign_lut_array := (
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
true, true, true, true, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false, 
false, false, false, false
);
constant EG_EG_DIFF_ETA_LUT_UFIXED : calo_calo_diff_eta_lut_ufixed_array := CALO_CALO_DIFF_ETA_LUT_UFIXED;
constant EG_TAU_DIFF_ETA_LUT_UFIXED : calo_calo_diff_eta_lut_ufixed_array := CALO_CALO_DIFF_ETA_LUT_UFIXED;
constant EG_JET_DIFF_ETA_LUT_UFIXED : calo_calo_diff_eta_lut_ufixed_array := CALO_CALO_DIFF_ETA_LUT_UFIXED;
constant JET_EG_DIFF_ETA_LUT_UFIXED : calo_calo_diff_eta_lut_ufixed_array := CALO_CALO_DIFF_ETA_LUT_UFIXED;
constant JET_JET_DIFF_ETA_LUT_UFIXED : calo_calo_diff_eta_lut_ufixed_array := CALO_CALO_DIFF_ETA_LUT_UFIXED;
constant JET_TAU_DIFF_ETA_LUT_UFIXED : calo_calo_diff_eta_lut_ufixed_array := CALO_CALO_DIFF_ETA_LUT_UFIXED;
constant TAU_EG_DIFF_ETA_LUT_UFIXED : calo_calo_diff_eta_lut_ufixed_array := CALO_CALO_DIFF_ETA_LUT_UFIXED;
constant TAU_JET_DIFF_ETA_LUT_UFIXED : calo_calo_diff_eta_lut_ufixed_array := CALO_CALO_DIFF_ETA_LUT_UFIXED;
constant TAU_TAU_DIFF_ETA_LUT_UFIXED : calo_calo_diff_eta_lut_ufixed_array := CALO_CALO_DIFF_ETA_LUT_UFIXED;
constant EG_EG_DIFF_PHI_LUT_UFIXED : calo_calo_diff_phi_lut_ufixed_array := CALO_CALO_DIFF_PHI_LUT_UFIXED;
constant EG_TAU_DIFF_PHI_LUT_UFIXED : calo_calo_diff_phi_lut_ufixed_array := CALO_CALO_DIFF_PHI_LUT_UFIXED;
constant EG_JET_DIFF_PHI_LUT_UFIXED : calo_calo_diff_phi_lut_ufixed_array := CALO_CALO_DIFF_PHI_LUT_UFIXED;
constant JET_EG_DIFF_PHI_LUT_UFIXED : calo_calo_diff_phi_lut_ufixed_array := CALO_CALO_DIFF_PHI_LUT_UFIXED;
constant JET_JET_DIFF_PHI_LUT_UFIXED : calo_calo_diff_phi_lut_ufixed_array := CALO_CALO_DIFF_PHI_LUT_UFIXED;
constant JET_TAU_DIFF_PHI_LUT_UFIXED : calo_calo_diff_phi_lut_ufixed_array := CALO_CALO_DIFF_PHI_LUT_UFIXED;
constant TAU_EG_DIFF_PHI_LUT_UFIXED : calo_calo_diff_phi_lut_ufixed_array := CALO_CALO_DIFF_PHI_LUT_UFIXED;
constant TAU_JET_DIFF_PHI_LUT_UFIXED : calo_calo_diff_phi_lut_ufixed_array := CALO_CALO_DIFF_PHI_LUT_UFIXED;
constant TAU_TAU_DIFF_PHI_LUT_UFIXED : calo_calo_diff_phi_lut_ufixed_array := CALO_CALO_DIFF_PHI_LUT_UFIXED;
constant TAU_PT_LUT_UFIXED : eg_pt_lut_ufixed_array := EG_PT_LUT_UFIXED;
constant EG_EG_COSH_DETA_LUT_UFIXED : calo_calo_cosh_deta_lut_ufixed_array := CALO_CALO_COSH_DETA_LUT_UFIXED;
constant EG_TAU_COSH_DETA_LUT_UFIXED : calo_calo_cosh_deta_lut_ufixed_array := CALO_CALO_COSH_DETA_LUT_UFIXED;
constant EG_JET_COSH_DETA_LUT_UFIXED : calo_calo_cosh_deta_lut_ufixed_array := CALO_CALO_COSH_DETA_LUT_UFIXED;
constant JET_EG_COSH_DETA_LUT_UFIXED : calo_calo_cosh_deta_lut_ufixed_array := CALO_CALO_COSH_DETA_LUT_UFIXED;
constant JET_JET_COSH_DETA_LUT_UFIXED : calo_calo_cosh_deta_lut_ufixed_array := CALO_CALO_COSH_DETA_LUT_UFIXED;
constant JET_TAU_COSH_DETA_LUT_UFIXED : calo_calo_cosh_deta_lut_ufixed_array := CALO_CALO_COSH_DETA_LUT_UFIXED;
constant TAU_EG_COSH_DETA_LUT_UFIXED : calo_calo_cosh_deta_lut_ufixed_array := CALO_CALO_COSH_DETA_LUT_UFIXED;
constant TAU_JET_COSH_DETA_LUT_UFIXED : calo_calo_cosh_deta_lut_ufixed_array := CALO_CALO_COSH_DETA_LUT_UFIXED;
constant TAU_TAU_COSH_DETA_LUT_UFIXED : calo_calo_cosh_deta_lut_ufixed_array := CALO_CALO_COSH_DETA_LUT_UFIXED;
constant EG_EG_COS_DPHI_LUT_UFIXED : calo_calo_cos_dphi_lut_ufixed_array := CALO_CALO_COS_DPHI_LUT_UFIXED;
constant EG_TAU_COS_DPHI_LUT_UFIXED : calo_calo_cos_dphi_lut_ufixed_array := CALO_CALO_COS_DPHI_LUT_UFIXED;
constant EG_JET_COS_DPHI_LUT_UFIXED : calo_calo_cos_dphi_lut_ufixed_array := CALO_CALO_COS_DPHI_LUT_UFIXED;
constant JET_EG_COS_DPHI_LUT_UFIXED : calo_calo_cos_dphi_lut_ufixed_array := CALO_CALO_COS_DPHI_LUT_UFIXED;
constant JET_JET_COS_DPHI_LUT_UFIXED : calo_calo_cos_dphi_lut_ufixed_array := CALO_CALO_COS_DPHI_LUT_UFIXED;
constant JET_TAU_COS_DPHI_LUT_UFIXED : calo_calo_cos_dphi_lut_ufixed_array := CALO_CALO_COS_DPHI_LUT_UFIXED;
constant TAU_EG_COS_DPHI_LUT_UFIXED : calo_calo_cos_dphi_lut_ufixed_array := CALO_CALO_COS_DPHI_LUT_UFIXED;
constant TAU_JET_COS_DPHI_LUT_UFIXED : calo_calo_cos_dphi_lut_ufixed_array := CALO_CALO_COS_DPHI_LUT_UFIXED;
constant TAU_TAU_COS_DPHI_LUT_UFIXED : calo_calo_cos_dphi_lut_ufixed_array := CALO_CALO_COS_DPHI_LUT_UFIXED;
constant EG_EG_COS_DPHI_SIGN_LUT : calo_calo_cos_dphi_sign_lut_array := CALO_CALO_COS_DPHI_SIGN_LUT;
constant EG_TAU_COS_DPHI_SIGN_LUT : calo_calo_cos_dphi_sign_lut_array := CALO_CALO_COS_DPHI_SIGN_LUT;
constant EG_JET_COS_DPHI_SIGN_LUT : calo_calo_cos_dphi_sign_lut_array := CALO_CALO_COS_DPHI_SIGN_LUT;
constant JET_EG_COS_DPHI_SIGN_LUT : calo_calo_cos_dphi_sign_lut_array := CALO_CALO_COS_DPHI_SIGN_LUT;
constant JET_JET_COS_DPHI_SIGN_LUT : calo_calo_cos_dphi_sign_lut_array := CALO_CALO_COS_DPHI_SIGN_LUT;
constant JET_TAU_COS_DPHI_SIGN_LUT : calo_calo_cos_dphi_sign_lut_array := CALO_CALO_COS_DPHI_SIGN_LUT;
constant TAU_EG_COS_DPHI_SIGN_LUT : calo_calo_cos_dphi_sign_lut_array := CALO_CALO_COS_DPHI_SIGN_LUT;
constant TAU_JET_COS_DPHI_SIGN_LUT : calo_calo_cos_dphi_sign_lut_array := CALO_CALO_COS_DPHI_SIGN_LUT;
constant TAU_TAU_COS_DPHI_SIGN_LUT : calo_calo_cos_dphi_sign_lut_array := CALO_CALO_COS_DPHI_SIGN_LUT;

end package;

