--------------------------------------------------------------------------------
-- Synthesizer : ISE 14.6
-- Platform    : Linux Ubuntu 10.04
-- Targets     : Synthese
--------------------------------------------------------------------------------
-- This work is held in copyright as an unpublished work by HEPHY (Institute
-- of High Energy Physics) All rights reserved.  This work may not be used
-- except by authorized licensees of HEPHY. This work is the
-- confidential information of HEPHY.
--------------------------------------------------------------------------------
-- $HeadURL: svn://heros.hephy.at/GlobalTriggerUpgrade/l1tm/L1Menu_CaloMuonCorrelation_2015_hb_test/vhdl/module_0/src/gtl_pkg.vhd $
-- $Date: 2015-08-24 11:49:40 +0200 (Mon, 24 Aug 2015) $
-- $Author: bergauer $
-- $Revision: 4173 $
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

use work.lhc_data_pkg.all;
use work.math_pkg.all;
-- use work.gt_mp7_core_pkg.all;
-- use work.l1tm_pkg.all;

package gtl_pkg is

-- Algorithms
constant NR_ALGOS : positive := 2; -- number of algorithmns (min. 32 for FDL registers width !!!) - written by TME
-- 
-- ==== FDL definitions - begin ============================================================
-- Definitions for prescalers (for FDL !)
-- constant PRESCALER_COUNTER_WIDTH : integer := 24;
-- type prescale_factor_array is array (NR_ALGOS-1 downto 0) of std_logic_vector(31 downto 0); -- same width as PCIe data
-- constant PRESCALE_FACTOR_INIT : ipb_regs_array(0 to MAX_NR_ALGOS-1) := ( others => X"00000001"); -- written by TME
-- 
-- -- Definitions for rate counters
-- constant RATE_COUNTER_WIDTH : integer := 32;
-- type rate_counter_array is array (NR_ALGOS-1 downto 0) of std_logic_vector(RATE_COUNTER_WIDTH-1 downto 0);
-- 
-- -- HB 2014-02-28: changed vector length of init values for finor- and veto-maks, because of min. 32 bits for register
-- constant MASKS_INIT : ipb_regs_array(0 to MAX_NR_ALGOS-1) := ( others => X"00000001"); --Finor and veto masks registers (bit 0 = finor, bit 1 = veto)
-- ==== FDL definitions - end ============================================================

-- ==== Versions - begin ============================================================
-- HB 2015-05-28: see l1tm_pkg.vhd in l1tm/...
-- constant L1TM_UID : std_logic_vector(127 downto 0) := X"00000000000000000000000000000000";
-- constant L1TM_NAME : std_logic_vector(128*8-1 downto 0) := X"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
-- constant L1TM_FW_UID : std_logic_vector(127 downto 0) := X"00000000000000000000000000000000";
-- 
-- -- Trigger Menu Editor software version - written by TME
-- constant L1TM_COMPILER_MAJOR_VERSION      : integer range 0 to 255 := 255;
-- constant L1TM_COMPILER_MINOR_VERSION      : integer range 0 to 255 := 255;
-- constant L1TM_COMPILER_REV_VERSION        : integer range 0 to 255 := 255;
-- constant L1TM_COMPILER_VERSION : std_logic_vector(31 downto 0) := X"00" &
--            std_logic_vector(to_unsigned(L1TM_COMPILER_MAJOR_VERSION, 8)) &
--            std_logic_vector(to_unsigned(L1TM_COMPILER_MINOR_VERSION, 8)) &
--            std_logic_vector(to_unsigned(L1TM_COMPILER_REV_VERSION, 8));
-- 
-- -- HB 2014-09-09: GTL and FDL firmware major, minor and revision versions moved to gt_mp7_core_pkg.vhd (GTL_FW_MAJOR_VERSION, etc.)
-- --                for creating a tag name by a script independent from L1Menu.
-- -- GTL firmware (fix part) version
-- constant GTL_FW_VERSION : std_logic_vector(31 downto 0) := X"00" &
--            std_logic_vector(to_unsigned(GTL_FW_MAJOR_VERSION, 8)) &
--            std_logic_vector(to_unsigned(GTL_FW_MINOR_VERSION, 8)) &
--            std_logic_vector(to_unsigned(GTL_FW_REV_VERSION, 8));
-- 
-- -- FDL firmware version
-- constant FDL_FW_VERSION : std_logic_vector(31 downto 0) := X"00" &
--            std_logic_vector(to_unsigned(FDL_FW_MAJOR_VERSION, 8)) &
--            std_logic_vector(to_unsigned(FDL_FW_MINOR_VERSION, 8)) &
--            std_logic_vector(to_unsigned(FDL_FW_REV_VERSION, 8));
-- 
-- ==== Versions - end ============================================================

-- ==== MUONs - begin ============================================================
-- MUONs
constant NR_MUON_TEMPLATES : positive range 1 to 4 := 4; -- number of max. templates for muon conditions
constant NR_MUON_OBJECTS : positive := MUON_ARRAY_LENGTH; -- from lhc_data_pkg.vhd
constant MAX_MUON_BITS : positive := MUON_DATA_WIDTH; -- from lhc_data_pkg.vhd

type d_s_i_muon_record is record
    charge_high, charge_low, iso_high, iso_low, eta_high, eta_low, qual_high, qual_low, pt_high, pt_low, phi_high, phi_low : natural range MAX_MUON_BITS-1 downto 0;
end record d_s_i_muon_record;

constant d_s_i_muon : d_s_i_muon_record := (35,34,33,32,31,23,22,19,18,10,9,0);

type muon_objects_array is array (natural range <>) of std_logic_vector(MAX_MUON_BITS-1 downto 0);
constant MAX_MUON_TEMPLATES_BITS : positive range 1 to MUON_DATA_WIDTH := 16;
type muon_templates_array is array (1 to NR_MUON_TEMPLATES) of std_logic_vector(MAX_MUON_TEMPLATES_BITS-1 downto 0);

-- type muon_templates_quality_array is array (1 to NR_MUON_TEMPLATES) of std_logic_vector((2**(d_s_i_muon.qual_high-d_s_i_muon.qual_low+1))-1 downto 0);
type muon_templates_quality_array is array (1 to NR_MUON_TEMPLATES) of std_logic_vector(15 downto 0);
-- type muon_templates_iso_array is array (1 to NR_MUON_TEMPLATES) of std_logic_vector((2**(d_s_i_muon.iso_high-d_s_i_muon.iso_low+1))-1 downto 0);
type muon_templates_iso_array is array (1 to NR_MUON_TEMPLATES) of std_logic_vector(3 downto 0);

type muon_templates_boolean_array is array (1 to NR_MUON_TEMPLATES) of boolean;
type muon_templates_string_array is array (1 to NR_MUON_TEMPLATES) of string(1 to 3);

-- HB 2014-04-15: types for muon_charge_correlations.vhd
type muon_charcorr_double_array is array (0 to NR_MUON_OBJECTS-1, 0 to NR_MUON_OBJECTS-1) of std_logic;
type muon_charcorr_triple_array is array (0 to NR_MUON_OBJECTS-1, 0 to NR_MUON_OBJECTS-1, 0 to NR_MUON_OBJECTS-1) of std_logic;
type muon_charcorr_quad_array is array (0 to NR_MUON_OBJECTS-1, 0 to NR_MUON_OBJECTS-1, 0 to NR_MUON_OBJECTS-1, 0 to NR_MUON_OBJECTS-1) of std_logic;
-- ==== MUONs - end ============================================================

-- ==== CALOs - begin ============================================================
-- CALOs
constant NR_CALO_TEMPLATES : positive range 1 to 4 := 4; -- number of max. templates for calorimeter conditions
constant NR_EG_OBJECTS : positive := EG_ARRAY_LENGTH; -- number eg objects, from lhc_data_pkg.vhd
constant NR_JET_OBJECTS : positive := JET_ARRAY_LENGTH; -- number jet objects, from lhc_data_pkg.vhd
constant NR_TAU_OBJECTS : positive := TAU_ARRAY_LENGTH; -- number tau objects, from lhc_data_pkg.vhd
constant MAX_CALO_BITS : positive := max(EG_DATA_WIDTH, JET_DATA_WIDTH, TAU_DATA_WIDTH);
constant MAX_ISO_BITS : positive range 1 to 2 := 2;

-- d_s_i_calo_record used for calo_conditions.vhd
type d_s_i_calo_record is record
    phi_high, phi_low, eta_high, eta_low, et_high, et_low : natural range MAX_CALO_BITS-1 downto 0;
end record d_s_i_calo_record;

constant d_s_i_eg : d_s_i_calo_record := (24,17,16,9,8,0);
constant d_s_i_jet : d_s_i_calo_record := (26,19,18,11,10,0);
constant d_s_i_tau : d_s_i_calo_record := (24,17,16,9,8,0);

-- HB 2015-02-16: changed for different "calo_records", each for eg, jet and tau.
-- different records used for calo_conditions_v2.vhd
-- used natural instead of string for object types
constant EG_TYPE : natural range 0 to 2 := 0;
constant JET_TYPE : natural range 0 to 2 := 1;
constant TAU_TYPE : natural range 0 to 2 := 2;

type d_s_i_eg_record is record
    iso_high, iso_low, phi_high, phi_low, eta_high, eta_low, et_high, et_low : natural range MAX_CALO_BITS-1 downto 0;
end record d_s_i_eg_record;

type d_s_i_jet_record is record
    phi_high, phi_low, eta_high, eta_low, et_high, et_low : natural range MAX_CALO_BITS-1 downto 0;
end record d_s_i_jet_record;

type d_s_i_tau_record is record
    iso_high, iso_low, phi_high, phi_low, eta_high, eta_low, et_high, et_low : natural range MAX_CALO_BITS-1 downto 0;
end record d_s_i_tau_record;

constant D_S_I_EG_V2: d_s_i_eg_record := (26,25,24,17,16,9,8,0);
constant D_S_I_JET_V2 : d_s_i_jet_record := (26,19,18,11,10,0);
constant D_S_I_TAU_V2 : d_s_i_tau_record := (26,25,24,17,16,9,8,0);

type calo_objects_array is array (natural range <>) of std_logic_vector(MAX_CALO_BITS-1 downto 0);
constant MAX_CALO_TEMPLATES_BITS : positive range 1 to MAX_CALO_BITS := 16;
type calo_templates_array is array (1 to NR_CALO_TEMPLATES) of std_logic_vector(MAX_CALO_TEMPLATES_BITS-1 downto 0);
type calo_templates_boolean_array is array (1 to NR_CALO_TEMPLATES) of boolean;
type calo_templates_iso_array is array (1 to NR_CALO_TEMPLATES) of std_logic_vector(2**MAX_ISO_BITS-1 downto 0);

-- ESUMs
constant MAX_ESUMS_BITS_TEMP : positive := max(ETT_DATA_WIDTH, HT_DATA_WIDTH, ETM_DATA_WIDTH);
constant MAX_ESUMS_BITS : positive := max(MAX_ESUMS_BITS_TEMP, HTM_DATA_WIDTH);
constant MAX_ESUMS_TEMPLATES_BITS : positive range 1 to MAX_ESUMS_BITS := 16;

constant ETT_TYPE : natural range 0 to 3 := 0;
constant HTT_TYPE : natural range 0 to 3 := 1;
constant ETM_TYPE : natural range 0 to 3 := 2;
constant HTM_TYPE : natural range 0 to 3 := 3;

type d_s_i_ett_record is record
    et_high, et_low : natural range MAX_ESUMS_BITS-1 downto 0;
end record d_s_i_ett_record;

type d_s_i_htt_record is record
    et_high, et_low : natural range MAX_ESUMS_BITS-1 downto 0;
end record d_s_i_htt_record;

type d_s_i_etm_record is record
    phi_high, phi_low, et_high, et_low : natural range MAX_ESUMS_BITS-1 downto 0;
end record d_s_i_etm_record;

type d_s_i_htm_record is record
    phi_high, phi_low, et_high, et_low : natural range MAX_ESUMS_BITS-1 downto 0;
end record d_s_i_htm_record;

constant D_S_I_ETT : d_s_i_ett_record := (11,0);
constant D_S_I_HTT : d_s_i_htt_record := (11,0);
constant D_S_I_ETM : d_s_i_etm_record := (19,12,11,0);
constant D_S_I_HTM : d_s_i_htm_record := (19,12,11,0);
-- ==== CALOs - end ============================================================
-- Correlations

-- Subtractors
constant MAX_DIFF_BITS : positive := 16;
type diff_inputs_array is array (natural range <>) of std_logic_vector(MAX_DIFF_BITS-1 downto 0);
type diff_integer_inputs_array is array (natural range <>) of integer;
type diff_2dim_integer_array is array (natural range <>, natural range <>) of integer;

-- "External conditions" (former "Technical Triggers" and "External Algorithms") definitions
constant NR_EXTERNAL_CONDITIONS : positive := EXTERNAL_CONDITIONS_DATA_WIDTH; -- number of "External conditions" inputs (proposed max. NR_EXTERNAL_CONDITIONS = 256), from lhc_data_pkg.vhd

-- Parameter for sub_eta_obj_vs_obj and sub_phi_obj_vs_obj instances of correlation conditions

constant PI : real :=  3.14159;

constant PHI_HALF_RANGE_REAL : real := PI;
constant ETA_RANGE_REAL : real := 10.0; -- eta range max.: -5.0 to +5.0
subtype dr_squared_range_real is real range 0.0 to ((ETA_RANGE_REAL**2)+(PHI_HALF_RANGE_REAL**2));
subtype diff_eta_range_real is real range -ETA_RANGE_REAL to ETA_RANGE_REAL;
subtype diff_phi_range_real is real range 0.0 to PHI_HALF_RANGE_REAL;

constant POSITION_FINAL_PRECISION : positive := 3; -- 3 => max. number, higher numbers exceed 32 bit integer values !!!

-- HB 2015-08-17: LUT for eta values (values are in the center of bins).
subtype eta_range_integer is integer range -5000 to 5000;

type eg_eta_lut_array is array (0 to 255) of eta_range_integer;
constant eg_eta_lut : eg_eta_lut_array := (
22, 66, 109, 153, 196, 240, 283, 327, 370, 414, 457, 501, 544, 588, 631, 675,
718, 762, 805, 849, 892, 936, 979, 1023, 1066, 1110, 1153, 1197, 1240, 1284, 1327, 1371,
1414, 1458, 1501, 1545, 1588, 1632, 1675, 1719, 1762, 1806, 1849, 1893, 1936, 1980, 2023, 2067,
2110, 2154, 2197, 2241, 2284, 2328, 2371, 2415, 2458, 2502, 2545, 2589, 2632, 2676, 2719, 2763,
2806, 2850, 2893, 2937, 2980, 3024, 3067, 3111, 3154, 3198, 3241, 3285, 3328, 3372, 3415, 3459,
3502, 3546, 3589, 3633, 3676, 3720, 3763, 3807, 3850, 3894, 3937, 3981, 4024, 4068, 4111, 4155,
4198, 4242, 4285, 4329, 4372, 4416, 4459, 4503, 4546, 4590, 4633, 4677, 4720, 4764, 4807, 4851,
4894, 4938, 4981, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -- eta range -5.0 to 5.0
0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4981, -4938, -4894,
-4851, -4807, -4764, -4720, -4677, -4633, -4590, -4546, -4503, -4459, -4416, -4372, -4329, -4285, -4242, -4198,
-4155, -4111, -4068, -4024, -3981, -3937, -3894, -3850, -3807, -3763, -3720, -3676, -3633, -3589, -3546, -3502,
-3459, -3415, -3372, -3328, -3285, -3241, -3198, -3154, -3111, -3067, -3024, -2980, -2937, -2893, -2850, -2806,
-2763, -2719, -2676, -2632, -2589, -2545, -2502, -2458, -2415, -2371, -2328, -2284, -2241, -2197, -2154, -2110,
-2067, -2023, -1980, -1936, -1893, -1849, -1806, -1762, -1719, -1675, -1632, -1588, -1545, -1501, -1458, -1414,
-1371, -1327, -1284, -1240, -1197, -1153, -1110, -1066, -1023, -979, -936, -892, -849, -805, -762, -718,
-675, -631, -588, -544, -501, -457, -414, -370, -327, -283, -240, -196, -153, -109, -66, -22
);

type tau_eta_lut_array is array (0 to 255) of eta_range_integer;
constant tau_eta_lut : tau_eta_lut_array := (
22, 66, 109, 153, 196, 240, 283, 327, 370, 414, 457, 501, 544, 588, 631, 675,
718, 762, 805, 849, 892, 936, 979, 1023, 1066, 1110, 1153, 1197, 1240, 1284, 1327, 1371,
1414, 1458, 1501, 1545, 1588, 1632, 1675, 1719, 1762, 1806, 1849, 1893, 1936, 1980, 2023, 2067,
2110, 2154, 2197, 2241, 2284, 2328, 2371, 2415, 2458, 2502, 2545, 2589, 2632, 2676, 2719, 2763,
2806, 2850, 2893, 2937, 2980, 3024, 3067, 3111, 3154, 3198, 3241, 3285, 3328, 3372, 3415, 3459,
3502, 3546, 3589, 3633, 3676, 3720, 3763, 3807, 3850, 3894, 3937, 3981, 4024, 4068, 4111, 4155,
4198, 4242, 4285, 4329, 4372, 4416, 4459, 4503, 4546, 4590, 4633, 4677, 4720, 4764, 4807, 4851,
4894, 4938, 4981, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -- eta range -5.0 to 5.0
0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4981, -4938, -4894,
-4851, -4807, -4764, -4720, -4677, -4633, -4590, -4546, -4503, -4459, -4416, -4372, -4329, -4285, -4242, -4198,
-4155, -4111, -4068, -4024, -3981, -3937, -3894, -3850, -3807, -3763, -3720, -3676, -3633, -3589, -3546, -3502,
-3459, -3415, -3372, -3328, -3285, -3241, -3198, -3154, -3111, -3067, -3024, -2980, -2937, -2893, -2850, -2806,
-2763, -2719, -2676, -2632, -2589, -2545, -2502, -2458, -2415, -2371, -2328, -2284, -2241, -2197, -2154, -2110,
-2067, -2023, -1980, -1936, -1893, -1849, -1806, -1762, -1719, -1675, -1632, -1588, -1545, -1501, -1458, -1414,
-1371, -1327, -1284, -1240, -1197, -1153, -1110, -1066, -1023, -979, -936, -892, -849, -805, -762, -718,
-675, -631, -588, -544, -501, -457, -414, -370, -327, -283, -240, -196, -153, -109, -66, -22
);

type muon_eta_lut_array is array (0 to 511) of eta_range_integer;
constant muon_eta_lut : muon_eta_lut_array := (
6, 17, 28, 39, 49, 60, 71, 82, 93, 104, 115, 126, 136, 147, 158, 169,
180, 191, 202, 213, 223, 234, 245, 256, 267, 278, 289, 300, 310, 321, 332, 343,
354, 365, 376, 387, 397, 408, 419, 430, 441, 452, 463, 474, 484, 495, 506, 517,
528, 539, 550, 561, 571, 582, 593, 604, 615, 626, 637, 648, 658, 669, 680, 691,
702, 713, 724, 735, 745, 756, 767, 778, 789, 800, 811, 822, 832, 843, 854, 865,
876, 887, 898, 909, 919, 930, 941, 952, 963, 974, 985, 996, 1006, 1017, 1028, 1039,
1050, 1061, 1072, 1083, 1093, 1104, 1115, 1126, 1137, 1148, 1159, 1170, 1180, 1191, 1202, 1213,
1224, 1235, 1246, 1257, 1267, 1278, 1289, 1300, 1311, 1322, 1333, 1344, 1354, 1365, 1376, 1387,
1398, 1409, 1420, 1431, 1441, 1452, 1463, 1474, 1485, 1496, 1507, 1518, 1528, 1539, 1550, 1561,
1572, 1583, 1594, 1605, 1615, 1626, 1637, 1648, 1659, 1670, 1681, 1692, 1702, 1713, 1724, 1735,
1746, 1757, 1768, 1779, 1789, 1800, 1811, 1822, 1833, 1844, 1855, 1866, 1876, 1887, 1898, 1909,
1920, 1931, 1942, 1953, 1963, 1974, 1985, 1996, 2007, 2018, 2029, 2040, 2050, 2061, 2072, 2083,
2094, 2105, 2116, 2127, 2137, 2148, 2159, 2170, 2181, 2192, 2203, 2214, 2224, 2235, 2246, 2257,
2268, 2279, 2290, 2301, 2311, 2322, 2333, 2344, 2355, 2366, 2377, 2388, 2398, 2409, 2420, 2431,
2442, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -- eta range -2.45 to 2.45
0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0, -2442,
-2431, -2420, -2409, -2398, -2388, -2377, -2366, -2355, -2344, -2333, -2322, -2311, -2301, -2290, -2279, -2268,
-2257, -2246, -2235, -2224, -2214, -2203, -2192, -2181, -2170, -2159, -2148, -2137, -2127, -2116, -2105, -2094,
-2083, -2072, -2061, -2050, -2040, -2029, -2018, -2007, -1996, -1985, -1974, -1963, -1953, -1942, -1931, -1920,
-1909, -1898, -1887, -1876, -1866, -1855, -1844, -1833, -1822, -1811, -1800, -1789, -1779, -1768, -1757, -1746,
-1735, -1724, -1713, -1702, -1692, -1681, -1670, -1659, -1648, -1637, -1626, -1615, -1605, -1594, -1583, -1572,
-1561, -1550, -1539, -1528, -1518, -1507, -1496, -1485, -1474, -1463, -1452, -1441, -1431, -1420, -1409, -1398,
-1387, -1376, -1365, -1354, -1344, -1333, -1322, -1311, -1300, -1289, -1278, -1267, -1257, -1246, -1235, -1224,
-1213, -1202, -1191, -1180, -1170, -1159, -1148, -1137, -1126, -1115, -1104, -1093, -1083, -1072, -1061, -1050,
-1039, -1028, -1017, -1006, -996, -985, -974, -963, -952, -941, -930, -919, -909, -898, -887, -876,
-865, -854, -843, -832, -822, -811, -800, -789, -778, -767, -756, -745, -735, -724, -713, -702,
-691, -680, -669, -658, -648, -637, -626, -615, -604, -593, -582, -571, -561, -550, -539, -528,
-517, -506, -495, -484, -474, -463, -452, -441, -430, -419, -408, -397, -387, -376, -365, -354,
-343, -332, -321, -310, -300, -289, -278, -267, -256, -245, -234, -223, -213, -202, -191, -180,
-169, -158, -147, -136, -126, -115, -104, -93, -82, -71, -60, -49, -39, -28, -17, -6
);

constant PHI_HALF_RANGE_INTEGER : positive := 3142; -- or 31415, depends on how many digits after comma used;
subtype phi_range_integer is natural range 0 to 6283;

-- HB 2015-08-17: LUT for eta values (values are in the center of bins).
type eg_phi_lut_array is array (0 to 255) of phi_range_integer;
constant eg_phi_lut : eg_phi_lut_array := (
22, 66, 110, 153, 197, 240, 284, 328, 371, 415, 459, 502, 546, 590, 633, 677,
720, 764, 808, 851, 895, 939, 982, 1026, 1070, 1113, 1157, 1200, 1244, 1288, 1331, 1375,
1419, 1462, 1506, 1549, 1593, 1637, 1680, 1724, 1768, 1811, 1855, 1899, 1942, 1986, 2029, 2073,
2117, 2160, 2204, 2248, 2291, 2335, 2379, 2422, 2466, 2509, 2553, 2597, 2640, 2684, 2728, 2771,
2815, 2858, 2902, 2946, 2989, 3033, 3077, 3120, 3164, 3208, 3251, 3295, 3338, 3382, 3426, 3469,
3513, 3557, 3600, 3644, 3688, 3731, 3775, 3818, 3862, 3906, 3949, 3993, 4037, 4080, 4124, 4167,
4211, 4255, 4298, 4342, 4386, 4429, 4473, 4517, 4560, 4604, 4647, 4691, 4735, 4778, 4822, 4866,
4909, 4953, 4997, 5040, 5084, 5127, 5171, 5215, 5258, 5302, 5346, 5389, 5433, 5476, 5520, 5564,
5607, 5651, 5695, 5738, 5782, 5826, 5869, 5913, 5956, 6000, 6044, 6087, 6131, 6175, 6218, 6262, -- phi range 0 to 2*PI=6.283
0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0
);

type tau_phi_lut_array is array (0 to 255) of phi_range_integer;
constant tau_phi_lut : tau_phi_lut_array := (
22, 66, 110, 153, 197, 240, 284, 328, 371, 415, 459, 502, 546, 590, 633, 677,
720, 764, 808, 851, 895, 939, 982, 1026, 1070, 1113, 1157, 1200, 1244, 1288, 1331, 1375,
1419, 1462, 1506, 1549, 1593, 1637, 1680, 1724, 1768, 1811, 1855, 1899, 1942, 1986, 2029, 2073,
2117, 2160, 2204, 2248, 2291, 2335, 2379, 2422, 2466, 2509, 2553, 2597, 2640, 2684, 2728, 2771,
2815, 2858, 2902, 2946, 2989, 3033, 3077, 3120, 3164, 3208, 3251, 3295, 3338, 3382, 3426, 3469,
3513, 3557, 3600, 3644, 3688, 3731, 3775, 3818, 3862, 3906, 3949, 3993, 4037, 4080, 4124, 4167,
4211, 4255, 4298, 4342, 4386, 4429, 4473, 4517, 4560, 4604, 4647, 4691, 4735, 4778, 4822, 4866,
4909, 4953, 4997, 5040, 5084, 5127, 5171, 5215, 5258, 5302, 5346, 5389, 5433, 5476, 5520, 5564,
5607, 5651, 5695, 5738, 5782, 5826, 5869, 5913, 5956, 6000, 6044, 6087, 6131, 6175, 6218, 6262,
0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -- phi range 0 to 2*PI=6.283
0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0
);

type muon_phi_lut_array is array (0 to 1023) of phi_range_integer;
constant muon_phi_lut : muon_phi_lut_array := (
6, 17, 28, 39, 50, 60, 71, 82, 93, 104, 115, 126, 137, 148, 159, 170,
180, 191, 202, 213, 224, 235, 246, 257, 268, 279, 290, 300, 311, 322, 333, 344,
355, 366, 377, 388, 399, 410, 420, 431, 442, 453, 464, 475, 486, 497, 508, 519,
530, 540, 551, 562, 573, 584, 595, 606, 617, 628, 639, 650, 660, 671, 682, 693,
704, 715, 726, 737, 748, 759, 770, 780, 791, 802, 813, 824, 835, 846, 857, 868,
879, 890, 900, 911, 922, 933, 944, 955, 966, 977, 988, 999, 1010, 1020, 1031, 1042,
1053, 1064, 1075, 1086, 1097, 1108, 1119, 1130, 1140, 1151, 1162, 1173, 1184, 1195, 1206, 1217,
1228, 1239, 1250, 1260, 1271, 1282, 1293, 1304, 1315, 1326, 1337, 1348, 1359, 1369, 1380, 1391,
1402, 1413, 1424, 1435, 1446, 1457, 1468, 1479, 1489, 1500, 1511, 1522, 1533, 1544, 1555, 1566,
1577, 1588, 1599, 1609, 1620, 1631, 1642, 1653, 1664, 1675, 1686, 1697, 1708, 1719, 1729, 1740,
1751, 1762, 1773, 1784, 1795, 1806, 1817, 1828, 1839, 1849, 1860, 1871, 1882, 1893, 1904, 1915,
1926, 1937, 1948, 1959, 1969, 1980, 1991, 2002, 2013, 2024, 2035, 2046, 2057, 2068, 2079, 2089,
2100, 2111, 2122, 2133, 2144, 2155, 2166, 2177, 2188, 2199, 2209, 2220, 2231, 2242, 2253, 2264,
2275, 2286, 2297, 2308, 2319, 2329, 2340, 2351, 2362, 2373, 2384, 2395, 2406, 2417, 2428, 2439,
2449, 2460, 2471, 2482, 2493, 2504, 2515, 2526, 2537, 2548, 2558, 2569, 2580, 2591, 2602, 2613,
2624, 2635, 2646, 2657, 2668, 2678, 2689, 2700, 2711, 2722, 2733, 2744, 2755, 2766, 2777, 2788,
2798, 2809, 2820, 2831, 2842, 2853, 2864, 2875, 2886, 2897, 2908, 2918, 2929, 2940, 2951, 2962,
2973, 2984, 2995, 3006, 3017, 3028, 3038, 3049, 3060, 3071, 3082, 3093, 3104, 3115, 3126, 3137,
3148, 3158, 3169, 3180, 3191, 3202, 3213, 3224, 3235, 3246, 3257, 3268, 3278, 3289, 3300, 3311,
3322, 3333, 3344, 3355, 3366, 3377, 3388, 3398, 3409, 3420, 3431, 3442, 3453, 3464, 3475, 3486,
3497, 3508, 3518, 3529, 3540, 3551, 3562, 3573, 3584, 3595, 3606, 3617, 3628, 3638, 3649, 3660,
3671, 3682, 3693, 3704, 3715, 3726, 3737, 3748, 3758, 3769, 3780, 3791, 3802, 3813, 3824, 3835,
3846, 3857, 3867, 3878, 3889, 3900, 3911, 3922, 3933, 3944, 3955, 3966, 3977, 3987, 3998, 4009,
4020, 4031, 4042, 4053, 4064, 4075, 4086, 4097, 4107, 4118, 4129, 4140, 4151, 4162, 4173, 4184,
4195, 4206, 4217, 4227, 4238, 4249, 4260, 4271, 4282, 4293, 4304, 4315, 4326, 4337, 4347, 4358,
4369, 4380, 4391, 4402, 4413, 4424, 4435, 4446, 4457, 4467, 4478, 4489, 4500, 4511, 4522, 4533,
4544, 4555, 4566, 4577, 4587, 4598, 4609, 4620, 4631, 4642, 4653, 4664, 4675, 4686, 4697, 4707,
4718, 4729, 4740, 4751, 4762, 4773, 4784, 4795, 4806, 4817, 4827, 4838, 4849, 4860, 4871, 4882,
4893, 4904, 4915, 4926, 4937, 4947, 4958, 4969, 4980, 4991, 5002, 5013, 5024, 5035, 5046, 5056,
5067, 5078, 5089, 5100, 5111, 5122, 5133, 5144, 5155, 5166, 5176, 5187, 5198, 5209, 5220, 5231,
5242, 5253, 5264, 5275, 5286, 5296, 5307, 5318, 5329, 5340, 5351, 5362, 5373, 5384, 5395, 5406,
5416, 5427, 5438, 5449, 5460, 5471, 5482, 5493, 5504, 5515, 5526, 5536, 5547, 5558, 5569, 5580,
5591, 5602, 5613, 5624, 5635, 5646, 5656, 5667, 5678, 5689, 5700, 5711, 5722, 5733, 5744, 5755,
5766, 5776, 5787, 5798, 5809, 5820, 5831, 5842, 5853, 5864, 5875, 5886, 5896, 5907, 5918, 5929,
5940, 5951, 5962, 5973, 5984, 5995, 6006, 6016, 6027, 6038, 6049, 6060, 6071, 6082, 6093, 6104,
6115, 6126, 6136, 6147, 6158, 6169, 6180, 6191, 6202, 6213, 6224, 6235, 6246, 6256, 6267, 6278, -- phi range 0 to 2*PI=6.283
0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0
);

constant INV_MASS_COSH_COS_PRECISION : positive := 3; -- 3 digits after decimal point (after roundimg to the 5th digit)
constant INV_MASS_PT_PRECISION : positive := 1; -- 1 digit after decimal point

subtype eg_et_range_integer is integer range 0 to 2555;

-- type eg_et_lut_array is array (0 to 511) of eg_et_range_integer;
type eg_et_lut_array is array (0 to 2**(D_S_I_EG_V2.et_high-D_S_I_EG_V2.et_low+1)-1) of eg_et_range_integer;
constant EG_ET_LUT: eg_et_lut_array := (
0, 5, 10, 15, 20, 25, 30, 35, 40, 45, 50, 55, 60, 65, 70, 75,
80, 85, 90, 95, 100, 105, 110, 115, 120, 125, 130, 135, 140, 145, 150, 155,
160, 165, 170, 175, 180, 185, 190, 195, 200, 205, 210, 215, 220, 225, 230, 235,
240, 245, 250, 255, 260, 265, 270, 275, 280, 285, 290, 295, 300, 305, 310, 315,
320, 325, 330, 335, 340, 345, 350, 355, 360, 365, 370, 375, 380, 385, 390, 395,
400, 405, 410, 415, 420, 425, 430, 435, 440, 445, 450, 455, 460, 465, 470, 475,
480, 485, 490, 495, 500, 505, 510, 515, 520, 525, 530, 535, 540, 545, 550, 555,
560, 565, 570, 575, 580, 585, 590, 595, 600, 605, 610, 615, 620, 625, 630, 635,
640, 645, 650, 655, 660, 665, 670, 675, 680, 685, 690, 695, 700, 705, 710, 715,
720, 725, 730, 735, 740, 745, 750, 755, 760, 765, 770, 775, 780, 785, 790, 795,
800, 805, 810, 815, 820, 825, 830, 835, 840, 845, 850, 855, 860, 865, 870, 875,
880, 885, 890, 895, 900, 905, 910, 915, 920, 925, 930, 935, 940, 945, 950, 955,
960, 965, 970, 975, 980, 985, 990, 995, 1000, 1005, 1010, 1015, 1020, 1025, 1030, 1035,
1040, 1045, 1050, 1055, 1060, 1065, 1070, 1075, 1080, 1085, 1090, 1095, 1100, 1105, 1110, 1115,
1120, 1125, 1130, 1135, 1140, 1145, 1150, 1155, 1160, 1165, 1170, 1175, 1180, 1185, 1190, 1195,
1200, 1205, 1210, 1215, 1220, 1225, 1230, 1235, 1240, 1245, 1250, 1255, 1260, 1265, 1270, 1275,
1280, 1285, 1290, 1295, 1300, 1305, 1310, 1315, 1320, 1325, 1330, 1335, 1340, 1345, 1350, 1355,
1360, 1365, 1370, 1375, 1380, 1385, 1390, 1395, 1400, 1405, 1410, 1415, 1420, 1425, 1430, 1435,
1440, 1445, 1450, 1455, 1460, 1465, 1470, 1475, 1480, 1485, 1490, 1495, 1500, 1505, 1510, 1515,
1520, 1525, 1530, 1535, 1540, 1545, 1550, 1555, 1560, 1565, 1570, 1575, 1580, 1585, 1590, 1595,
1600, 1605, 1610, 1615, 1620, 1625, 1630, 1635, 1640, 1645, 1650, 1655, 1660, 1665, 1670, 1675,
1680, 1685, 1690, 1695, 1700, 1705, 1710, 1715, 1720, 1725, 1730, 1735, 1740, 1745, 1750, 1755,
1760, 1765, 1770, 1775, 1780, 1785, 1790, 1795, 1800, 1805, 1810, 1815, 1820, 1825, 1830, 1835,
1840, 1845, 1850, 1855, 1860, 1865, 1870, 1875, 1880, 1885, 1890, 1895, 1900, 1905, 1910, 1915,
1920, 1925, 1930, 1935, 1940, 1945, 1950, 1955, 1960, 1965, 1970, 1975, 1980, 1985, 1990, 1995,
2000, 2005, 2010, 2015, 2020, 2025, 2030, 2035, 2040, 2045, 2050, 2055, 2060, 2065, 2070, 2075,
2080, 2085, 2090, 2095, 2100, 2105, 2110, 2115, 2120, 2125, 2130, 2135, 2140, 2145, 2150, 2155,
2160, 2165, 2170, 2175, 2180, 2185, 2190, 2195, 2200, 2205, 2210, 2215, 2220, 2225, 2230, 2235,
2240, 2245, 2250, 2255, 2260, 2265, 2270, 2275, 2280, 2285, 2290, 2295, 2300, 2305, 2310, 2315,
2320, 2325, 2330, 2335, 2340, 2345, 2350, 2355, 2360, 2365, 2370, 2375, 2380, 2385, 2390, 2395,
2400, 2405, 2410, 2415, 2420, 2425, 2430, 2435, 2440, 2445, 2450, 2455, 2460, 2465, 2470, 2475,
2480, 2485, 2490, 2495, 2500, 2505, 2510, 2515, 2520, 2525, 2530, 2535, 2540, 2545, 2550, 2555
);

type calo_calo_cosh_deta_lut_array is array (0 to 255, 0 to 255) of integer;
constant CALO_CALO_COSH_DETA_LUT: calo_calo_cosh_deta_lut_array := (

(1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001),
(1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004),
(1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009),
(1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015),
(1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024),
(1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034),
(1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047),
(1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061),
(1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078),
(1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096),
(1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117),
(1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139),
(1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164),
(1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191),
(1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221),
(1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252),
(1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286),
(1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323),
(1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361),
(1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403),
(1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447),
(1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494),
(1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544),
(1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596),
(1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652),
(1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711),
(1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773),
(1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838),
(1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907),
(1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979),
(1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056),
(2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136),
(2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220),
(2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308),
(2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401),
(2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498),
(2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600),
(2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707),
(2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819),
(2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936),
(2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059),
(3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188),
(3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323),
(3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464),
(3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611),
(3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766),
(3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927),
(3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096),
(4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273),
(4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458),
(4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651),
(4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853),
(4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064),
(5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285),
(5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516),
(5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757),
(5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010),
(6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273),
(6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548),
(6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836),
(6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137),
(7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451),
(7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780),
(7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123),
(8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481),
(8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856),
(8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247),
(9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656),
(9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083),
(10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529),
(10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995),
(10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482),
(11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990),
(11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522),
(12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077),
(13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656),
(13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 3571900, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262),
(14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 3730706, 3571900, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894),
(14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 3896573, 3730706, 3571900, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555),
(15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4069815, 3896573, 3730706, 3571900, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245),
(16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4250759, 4069815, 3896573, 3730706, 3571900, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966),
(16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 4439748, 4250759, 4069815, 3896573, 3730706, 3571900, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719),
(17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 4637139, 4439748, 4250759, 4069815, 3896573, 3730706, 3571900, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506),
(18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 4843306, 4637139, 4439748, 4250759, 4069815, 3896573, 3730706, 3571900, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327),
(19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 5058639, 4843306, 4637139, 4439748, 4250759, 4069815, 3896573, 3730706, 3571900, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186),
(20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 5283546, 5058639, 4843306, 4637139, 4439748, 4250759, 4069815, 3896573, 3730706, 3571900, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082),
(21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 5518453, 5283546, 5058639, 4843306, 4637139, 4439748, 4250759, 4069815, 3896573, 3730706, 3571900, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018),
(22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 5763803, 5518453, 5283546, 5058639, 4843306, 4637139, 4439748, 4250759, 4069815, 3896573, 3730706, 3571900, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996),
(22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 6020062, 5763803, 5518453, 5283546, 5058639, 4843306, 4637139, 4439748, 4250759, 4069815, 3896573, 3730706, 3571900, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018),
(24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 6287714, 6020062, 5763803, 5518453, 5283546, 5058639, 4843306, 4637139, 4439748, 4250759, 4069815, 3896573, 3730706, 3571900, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085),
(25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 6567266, 6287714, 6020062, 5763803, 5518453, 5283546, 5058639, 4843306, 4637139, 4439748, 4250759, 4069815, 3896573, 3730706, 3571900, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199),
(26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 6859246, 6567266, 6287714, 6020062, 5763803, 5518453, 5283546, 5058639, 4843306, 4637139, 4439748, 4250759, 4069815, 3896573, 3730706, 3571900, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363),
(27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 7164208, 6859246, 6567266, 6287714, 6020062, 5763803, 5518453, 5283546, 5058639, 4843306, 4637139, 4439748, 4250759, 4069815, 3896573, 3730706, 3571900, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579),
(28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 7482729, 7164208, 6859246, 6567266, 6287714, 6020062, 5763803, 5518453, 5283546, 5058639, 4843306, 4637139, 4439748, 4250759, 4069815, 3896573, 3730706, 3571900, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848),
(29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 7815411, 7482729, 7164208, 6859246, 6567266, 6287714, 6020062, 5763803, 5518453, 5283546, 5058639, 4843306, 4637139, 4439748, 4250759, 4069815, 3896573, 3730706, 3571900, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175),
(31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 8162884, 7815411, 7482729, 7164208, 6859246, 6567266, 6287714, 6020062, 5763803, 5518453, 5283546, 5058639, 4843306, 4637139, 4439748, 4250759, 4069815, 3896573, 3730706, 3571900, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560),
(32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 8525806, 8162884, 7815411, 7482729, 7164208, 6859246, 6567266, 6287714, 6020062, 5763803, 5518453, 5283546, 5058639, 4843306, 4637139, 4439748, 4250759, 4069815, 3896573, 3730706, 3571900, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007),
(34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 8904863, 8525806, 8162884, 7815411, 7482729, 7164208, 6859246, 6567266, 6287714, 6020062, 5763803, 5518453, 5283546, 5058639, 4843306, 4637139, 4439748, 4250759, 4069815, 3896573, 3730706, 3571900, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518),
(35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 9300773, 8904863, 8525806, 8162884, 7815411, 7482729, 7164208, 6859246, 6567266, 6287714, 6020062, 5763803, 5518453, 5283546, 5058639, 4843306, 4637139, 4439748, 4250759, 4069815, 3896573, 3730706, 3571900, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097),
(37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 9714286, 9300773, 8904863, 8525806, 8162884, 7815411, 7482729, 7164208, 6859246, 6567266, 6287714, 6020062, 5763803, 5518453, 5283546, 5058639, 4843306, 4637139, 4439748, 4250759, 4069815, 3896573, 3730706, 3571900, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746),
(38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 10146183, 9714286, 9300773, 8904863, 8525806, 8162884, 7815411, 7482729, 7164208, 6859246, 6567266, 6287714, 6020062, 5763803, 5518453, 5283546, 5058639, 4843306, 4637139, 4439748, 4250759, 4069815, 3896573, 3730706, 3571900, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468),
(40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 10597282, 10146183, 9714286, 9300773, 8904863, 8525806, 8162884, 7815411, 7482729, 7164208, 6859246, 6567266, 6287714, 6020062, 5763803, 5518453, 5283546, 5058639, 4843306, 4637139, 4439748, 4250759, 4069815, 3896573, 3730706, 3571900, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266),
(42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 11068437, 10597282, 10146183, 9714286, 9300773, 8904863, 8525806, 8162884, 7815411, 7482729, 7164208, 6859246, 6567266, 6287714, 6020062, 5763803, 5518453, 5283546, 5058639, 4843306, 4637139, 4439748, 4250759, 4069815, 3896573, 3730706, 3571900, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145),
(44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 11560540, 11068437, 10597282, 10146183, 9714286, 9300773, 8904863, 8525806, 8162884, 7815411, 7482729, 7164208, 6859246, 6567266, 6287714, 6020062, 5763803, 5518453, 5283546, 5058639, 4843306, 4637139, 4439748, 4250759, 4069815, 3896573, 3730706, 3571900, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107),
(46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 12074521, 11560540, 11068437, 10597282, 10146183, 9714286, 9300773, 8904863, 8525806, 8162884, 7815411, 7482729, 7164208, 6859246, 6567266, 6287714, 6020062, 5763803, 5518453, 5283546, 5058639, 4843306, 4637139, 4439748, 4250759, 4069815, 3896573, 3730706, 3571900, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157),
(48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 12611354, 12074521, 11560540, 11068437, 10597282, 10146183, 9714286, 9300773, 8904863, 8525806, 8162884, 7815411, 7482729, 7164208, 6859246, 6567266, 6287714, 6020062, 5763803, 5518453, 5283546, 5058639, 4843306, 4637139, 4439748, 4250759, 4069815, 3896573, 3730706, 3571900, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297),
(50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 13172055, 12611354, 12074521, 11560540, 11068437, 10597282, 10146183, 9714286, 9300773, 8904863, 8525806, 8162884, 7815411, 7482729, 7164208, 6859246, 6567266, 6287714, 6020062, 5763803, 5518453, 5283546, 5058639, 4843306, 4637139, 4439748, 4250759, 4069815, 3896573, 3730706, 3571900, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533),
(52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 13757685, 13172055, 12611354, 12074521, 11560540, 11068437, 10597282, 10146183, 9714286, 9300773, 8904863, 8525806, 8162884, 7815411, 7482729, 7164208, 6859246, 6567266, 6287714, 6020062, 5763803, 5518453, 5283546, 5058639, 4843306, 4637139, 4439748, 4250759, 4069815, 3896573, 3730706, 3571900, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868),
(54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 14369351, 13757685, 13172055, 12611354, 12074521, 11560540, 11068437, 10597282, 10146183, 9714286, 9300773, 8904863, 8525806, 8162884, 7815411, 7482729, 7164208, 6859246, 6567266, 6287714, 6020062, 5763803, 5518453, 5283546, 5058639, 4843306, 4637139, 4439748, 4250759, 4069815, 3896573, 3730706, 3571900, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307),
(57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 15008212, 14369351, 13757685, 13172055, 12611354, 12074521, 11560540, 11068437, 10597282, 10146183, 9714286, 9300773, 8904863, 8525806, 8162884, 7815411, 7482729, 7164208, 6859246, 6567266, 6287714, 6020062, 5763803, 5518453, 5283546, 5058639, 4843306, 4637139, 4439748, 4250759, 4069815, 3896573, 3730706, 3571900, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855),
(59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 15675477, 15008212, 14369351, 13757685, 13172055, 12611354, 12074521, 11560540, 11068437, 10597282, 10146183, 9714286, 9300773, 8904863, 8525806, 8162884, 7815411, 7482729, 7164208, 6859246, 6567266, 6287714, 6020062, 5763803, 5518453, 5283546, 5058639, 4843306, 4637139, 4439748, 4250759, 4069815, 3896573, 3730706, 3571900, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516),
(62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 16372409, 15675477, 15008212, 14369351, 13757685, 13172055, 12611354, 12074521, 11560540, 11068437, 10597282, 10146183, 9714286, 9300773, 8904863, 8525806, 8162884, 7815411, 7482729, 7164208, 6859246, 6567266, 6287714, 6020062, 5763803, 5518453, 5283546, 5058639, 4843306, 4637139, 4439748, 4250759, 4069815, 3896573, 3730706, 3571900, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295),
(65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 17100326, 16372409, 15675477, 15008212, 14369351, 13757685, 13172055, 12611354, 12074521, 11560540, 11068437, 10597282, 10146183, 9714286, 9300773, 8904863, 8525806, 8162884, 7815411, 7482729, 7164208, 6859246, 6567266, 6287714, 6020062, 5763803, 5518453, 5283546, 5058639, 4843306, 4637139, 4439748, 4250759, 4069815, 3896573, 3730706, 3571900, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197),
(68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 17860607, 17100326, 16372409, 15675477, 15008212, 14369351, 13757685, 13172055, 12611354, 12074521, 11560540, 11068437, 10597282, 10146183, 9714286, 9300773, 8904863, 8525806, 8162884, 7815411, 7482729, 7164208, 6859246, 6567266, 6287714, 6020062, 5763803, 5518453, 5283546, 5058639, 4843306, 4637139, 4439748, 4250759, 4069815, 3896573, 3730706, 3571900, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229),
(71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 18654689, 17860607, 17100326, 16372409, 15675477, 15008212, 14369351, 13757685, 13172055, 12611354, 12074521, 11560540, 11068437, 10597282, 10146183, 9714286, 9300773, 8904863, 8525806, 8162884, 7815411, 7482729, 7164208, 6859246, 6567266, 6287714, 6020062, 5763803, 5518453, 5283546, 5058639, 4843306, 4637139, 4439748, 4250759, 4069815, 3896573, 3730706, 3571900, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396),
(74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 19484076, 18654689, 17860607, 17100326, 16372409, 15675477, 15008212, 14369351, 13757685, 13172055, 12611354, 12074521, 11560540, 11068437, 10597282, 10146183, 9714286, 9300773, 8904863, 8525806, 8162884, 7815411, 7482729, 7164208, 6859246, 6567266, 6287714, 6020062, 5763803, 5518453, 5283546, 5058639, 4843306, 4637139, 4439748, 4250759, 4069815, 3896573, 3730706, 3571900, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703),
(77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 20350338, 19484076, 18654689, 17860607, 17100326, 16372409, 15675477, 15008212, 14369351, 13757685, 13172055, 12611354, 12074521, 11560540, 11068437, 10597282, 10146183, 9714286, 9300773, 8904863, 8525806, 8162884, 7815411, 7482729, 7164208, 6859246, 6567266, 6287714, 6020062, 5763803, 5518453, 5283546, 5058639, 4843306, 4637139, 4439748, 4250759, 4069815, 3896573, 3730706, 3571900, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157),
(81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 21255114, 20350338, 19484076, 18654689, 17860607, 17100326, 16372409, 15675477, 15008212, 14369351, 13757685, 13172055, 12611354, 12074521, 11560540, 11068437, 10597282, 10146183, 9714286, 9300773, 8904863, 8525806, 8162884, 7815411, 7482729, 7164208, 6859246, 6567266, 6287714, 6020062, 5763803, 5518453, 5283546, 5058639, 4843306, 4637139, 4439748, 4250759, 4069815, 3896573, 3730706, 3571900, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765),
(84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 22200117, 21255114, 20350338, 19484076, 18654689, 17860607, 17100326, 16372409, 15675477, 15008212, 14369351, 13757685, 13172055, 12611354, 12074521, 11560540, 11068437, 10597282, 10146183, 9714286, 9300773, 8904863, 8525806, 8162884, 7815411, 7482729, 7164208, 6859246, 6567266, 6287714, 6020062, 5763803, 5518453, 5283546, 5058639, 4843306, 4637139, 4439748, 4250759, 4069815, 3896573, 3730706, 3571900, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534),
(88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 23187134, 22200117, 21255114, 20350338, 19484076, 18654689, 17860607, 17100326, 16372409, 15675477, 15008212, 14369351, 13757685, 13172055, 12611354, 12074521, 11560540, 11068437, 10597282, 10146183, 9714286, 9300773, 8904863, 8525806, 8162884, 7815411, 7482729, 7164208, 6859246, 6567266, 6287714, 6020062, 5763803, 5518453, 5283546, 5058639, 4843306, 4637139, 4439748, 4250759, 4069815, 3896573, 3730706, 3571900, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470),
(92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 24218033, 23187134, 22200117, 21255114, 20350338, 19484076, 18654689, 17860607, 17100326, 16372409, 15675477, 15008212, 14369351, 13757685, 13172055, 12611354, 12074521, 11560540, 11068437, 10597282, 10146183, 9714286, 9300773, 8904863, 8525806, 8162884, 7815411, 7482729, 7164208, 6859246, 6567266, 6287714, 6020062, 5763803, 5518453, 5283546, 5058639, 4843306, 4637139, 4439748, 4250759, 4069815, 3896573, 3730706, 3571900, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581),
(96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 25294767, 24218033, 23187134, 22200117, 21255114, 20350338, 19484076, 18654689, 17860607, 17100326, 16372409, 15675477, 15008212, 14369351, 13757685, 13172055, 12611354, 12074521, 11560540, 11068437, 10597282, 10146183, 9714286, 9300773, 8904863, 8525806, 8162884, 7815411, 7482729, 7164208, 6859246, 6567266, 6287714, 6020062, 5763803, 5518453, 5283546, 5058639, 4843306, 4637139, 4439748, 4250759, 4069815, 3896573, 3730706, 3571900, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359, 100875),
(100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 26419372, 25294767, 24218033, 23187134, 22200117, 21255114, 20350338, 19484076, 18654689, 17860607, 17100326, 16372409, 15675477, 15008212, 14369351, 13757685, 13172055, 12611354, 12074521, 11560540, 11068437, 10597282, 10146183, 9714286, 9300773, 8904863, 8525806, 8162884, 7815411, 7482729, 7164208, 6859246, 6567266, 6287714, 6020062, 5763803, 5518453, 5283546, 5058639, 4843306, 4637139, 4439748, 4250759, 4069815, 3896573, 3730706, 3571900, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043, 105359),
(105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 27593977, 26419372, 25294767, 24218033, 23187134, 22200117, 21255114, 20350338, 19484076, 18654689, 17860607, 17100326, 16372409, 15675477, 15008212, 14369351, 13757685, 13172055, 12611354, 12074521, 11560540, 11068437, 10597282, 10146183, 9714286, 9300773, 8904863, 8525806, 8162884, 7815411, 7482729, 7164208, 6859246, 6567266, 6287714, 6020062, 5763803, 5518453, 5283546, 5058639, 4843306, 4637139, 4439748, 4250759, 4069815, 3896573, 3730706, 3571900, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936, 110043),
(110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 28820806, 27593977, 26419372, 25294767, 24218033, 23187134, 22200117, 21255114, 20350338, 19484076, 18654689, 17860607, 17100326, 16372409, 15675477, 15008212, 14369351, 13757685, 13172055, 12611354, 12074521, 11560540, 11068437, 10597282, 10146183, 9714286, 9300773, 8904863, 8525806, 8162884, 7815411, 7482729, 7164208, 6859246, 6567266, 6287714, 6020062, 5763803, 5518453, 5283546, 5058639, 4843306, 4637139, 4439748, 4250759, 4069815, 3896573, 3730706, 3571900, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045, 114936),
(114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 30102178, 28820806, 27593977, 26419372, 25294767, 24218033, 23187134, 22200117, 21255114, 20350338, 19484076, 18654689, 17860607, 17100326, 16372409, 15675477, 15008212, 14369351, 13757685, 13172055, 12611354, 12074521, 11560540, 11068437, 10597282, 10146183, 9714286, 9300773, 8904863, 8525806, 8162884, 7815411, 7482729, 7164208, 6859246, 6567266, 6287714, 6020062, 5763803, 5518453, 5283546, 5058639, 4843306, 4637139, 4439748, 4250759, 4069815, 3896573, 3730706, 3571900, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382, 120045),
(120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 31440521, 30102178, 28820806, 27593977, 26419372, 25294767, 24218033, 23187134, 22200117, 21255114, 20350338, 19484076, 18654689, 17860607, 17100326, 16372409, 15675477, 15008212, 14369351, 13757685, 13172055, 12611354, 12074521, 11560540, 11068437, 10597282, 10146183, 9714286, 9300773, 8904863, 8525806, 8162884, 7815411, 7482729, 7164208, 6859246, 6567266, 6287714, 6020062, 5763803, 5518453, 5283546, 5058639, 4843306, 4637139, 4439748, 4250759, 4069815, 3896573, 3730706, 3571900, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957, 125382),
(125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 32838366, 31440521, 30102178, 28820806, 27593977, 26419372, 25294767, 24218033, 23187134, 22200117, 21255114, 20350338, 19484076, 18654689, 17860607, 17100326, 16372409, 15675477, 15008212, 14369351, 13757685, 13172055, 12611354, 12074521, 11560540, 11068437, 10597282, 10146183, 9714286, 9300773, 8904863, 8525806, 8162884, 7815411, 7482729, 7164208, 6859246, 6567266, 6287714, 6020062, 5763803, 5518453, 5283546, 5058639, 4843306, 4637139, 4439748, 4250759, 4069815, 3896573, 3730706, 3571900, 3419853, 3274279, 3134901, 3001456, 2873692, 2751366, 2634248, 2522114, 2414754, 2311964, 2213550, 2119325, 2029111, 1942737, 1860039, 1780862, 1705055, 1632476, 1562985, 1496453, 1432753, 1371764, 1313372, 1257465, 1203938, 1152689, 1103622, 1056644, 1011665, 968601, 927370, 887895, 850099, 813913, 779267, 746095, 714336, 683928, 654815, 626942, 600254, 574703, 550240, 526817, 504392, 482921, 462365, 442683, 423839, 405798, 388524, 371985, 356151, 340991, 326476, 312578, 299273, 286534, 274337, 262659, 251478, 240774, 230525, 220712, 211317, 202322, 193709, 185464, 177569, 170011, 162774, 155845, 149211, 142860, 136779, 130957),
(130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 3571900, 3730706, 3896573, 4069815, 4250759, 4439748, 4637139, 4843306, 5058639, 5283546, 5518453, 5763803, 6020062, 6287714, 6567266, 6859246, 7164208, 7482729, 7815411, 8162884, 8525806, 8904863, 9300773, 9714286, 10146183, 10597282, 11068437, 11560540, 12074521, 12611354, 13172055, 13757685, 14369351, 15008212, 15675477, 16372409, 17100326, 17860607, 18654689, 19484076, 20350338, 21255114, 22200117, 23187134, 24218033, 25294767, 26419372, 27593977, 28820806, 30102178, 31440521, 32838366, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382),
(125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 3571900, 3730706, 3896573, 4069815, 4250759, 4439748, 4637139, 4843306, 5058639, 5283546, 5518453, 5763803, 6020062, 6287714, 6567266, 6859246, 7164208, 7482729, 7815411, 8162884, 8525806, 8904863, 9300773, 9714286, 10146183, 10597282, 11068437, 11560540, 12074521, 12611354, 13172055, 13757685, 14369351, 15008212, 15675477, 16372409, 17100326, 17860607, 18654689, 19484076, 20350338, 21255114, 22200117, 23187134, 24218033, 25294767, 26419372, 27593977, 28820806, 30102178, 31440521, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045),
(120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 3571900, 3730706, 3896573, 4069815, 4250759, 4439748, 4637139, 4843306, 5058639, 5283546, 5518453, 5763803, 6020062, 6287714, 6567266, 6859246, 7164208, 7482729, 7815411, 8162884, 8525806, 8904863, 9300773, 9714286, 10146183, 10597282, 11068437, 11560540, 12074521, 12611354, 13172055, 13757685, 14369351, 15008212, 15675477, 16372409, 17100326, 17860607, 18654689, 19484076, 20350338, 21255114, 22200117, 23187134, 24218033, 25294767, 26419372, 27593977, 28820806, 30102178, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936),
(114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 3571900, 3730706, 3896573, 4069815, 4250759, 4439748, 4637139, 4843306, 5058639, 5283546, 5518453, 5763803, 6020062, 6287714, 6567266, 6859246, 7164208, 7482729, 7815411, 8162884, 8525806, 8904863, 9300773, 9714286, 10146183, 10597282, 11068437, 11560540, 12074521, 12611354, 13172055, 13757685, 14369351, 15008212, 15675477, 16372409, 17100326, 17860607, 18654689, 19484076, 20350338, 21255114, 22200117, 23187134, 24218033, 25294767, 26419372, 27593977, 28820806, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043),
(110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 3571900, 3730706, 3896573, 4069815, 4250759, 4439748, 4637139, 4843306, 5058639, 5283546, 5518453, 5763803, 6020062, 6287714, 6567266, 6859246, 7164208, 7482729, 7815411, 8162884, 8525806, 8904863, 9300773, 9714286, 10146183, 10597282, 11068437, 11560540, 12074521, 12611354, 13172055, 13757685, 14369351, 15008212, 15675477, 16372409, 17100326, 17860607, 18654689, 19484076, 20350338, 21255114, 22200117, 23187134, 24218033, 25294767, 26419372, 27593977, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359),
(105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 3571900, 3730706, 3896573, 4069815, 4250759, 4439748, 4637139, 4843306, 5058639, 5283546, 5518453, 5763803, 6020062, 6287714, 6567266, 6859246, 7164208, 7482729, 7815411, 8162884, 8525806, 8904863, 9300773, 9714286, 10146183, 10597282, 11068437, 11560540, 12074521, 12611354, 13172055, 13757685, 14369351, 15008212, 15675477, 16372409, 17100326, 17860607, 18654689, 19484076, 20350338, 21255114, 22200117, 23187134, 24218033, 25294767, 26419372, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875),
(100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 3571900, 3730706, 3896573, 4069815, 4250759, 4439748, 4637139, 4843306, 5058639, 5283546, 5518453, 5763803, 6020062, 6287714, 6567266, 6859246, 7164208, 7482729, 7815411, 8162884, 8525806, 8904863, 9300773, 9714286, 10146183, 10597282, 11068437, 11560540, 12074521, 12611354, 13172055, 13757685, 14369351, 15008212, 15675477, 16372409, 17100326, 17860607, 18654689, 19484076, 20350338, 21255114, 22200117, 23187134, 24218033, 25294767, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581),
(96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 3571900, 3730706, 3896573, 4069815, 4250759, 4439748, 4637139, 4843306, 5058639, 5283546, 5518453, 5763803, 6020062, 6287714, 6567266, 6859246, 7164208, 7482729, 7815411, 8162884, 8525806, 8904863, 9300773, 9714286, 10146183, 10597282, 11068437, 11560540, 12074521, 12611354, 13172055, 13757685, 14369351, 15008212, 15675477, 16372409, 17100326, 17860607, 18654689, 19484076, 20350338, 21255114, 22200117, 23187134, 24218033, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470),
(92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 3571900, 3730706, 3896573, 4069815, 4250759, 4439748, 4637139, 4843306, 5058639, 5283546, 5518453, 5763803, 6020062, 6287714, 6567266, 6859246, 7164208, 7482729, 7815411, 8162884, 8525806, 8904863, 9300773, 9714286, 10146183, 10597282, 11068437, 11560540, 12074521, 12611354, 13172055, 13757685, 14369351, 15008212, 15675477, 16372409, 17100326, 17860607, 18654689, 19484076, 20350338, 21255114, 22200117, 23187134, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534),
(88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 3571900, 3730706, 3896573, 4069815, 4250759, 4439748, 4637139, 4843306, 5058639, 5283546, 5518453, 5763803, 6020062, 6287714, 6567266, 6859246, 7164208, 7482729, 7815411, 8162884, 8525806, 8904863, 9300773, 9714286, 10146183, 10597282, 11068437, 11560540, 12074521, 12611354, 13172055, 13757685, 14369351, 15008212, 15675477, 16372409, 17100326, 17860607, 18654689, 19484076, 20350338, 21255114, 22200117, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765),
(84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 3571900, 3730706, 3896573, 4069815, 4250759, 4439748, 4637139, 4843306, 5058639, 5283546, 5518453, 5763803, 6020062, 6287714, 6567266, 6859246, 7164208, 7482729, 7815411, 8162884, 8525806, 8904863, 9300773, 9714286, 10146183, 10597282, 11068437, 11560540, 12074521, 12611354, 13172055, 13757685, 14369351, 15008212, 15675477, 16372409, 17100326, 17860607, 18654689, 19484076, 20350338, 21255114, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157),
(81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 3571900, 3730706, 3896573, 4069815, 4250759, 4439748, 4637139, 4843306, 5058639, 5283546, 5518453, 5763803, 6020062, 6287714, 6567266, 6859246, 7164208, 7482729, 7815411, 8162884, 8525806, 8904863, 9300773, 9714286, 10146183, 10597282, 11068437, 11560540, 12074521, 12611354, 13172055, 13757685, 14369351, 15008212, 15675477, 16372409, 17100326, 17860607, 18654689, 19484076, 20350338, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703),
(77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 3571900, 3730706, 3896573, 4069815, 4250759, 4439748, 4637139, 4843306, 5058639, 5283546, 5518453, 5763803, 6020062, 6287714, 6567266, 6859246, 7164208, 7482729, 7815411, 8162884, 8525806, 8904863, 9300773, 9714286, 10146183, 10597282, 11068437, 11560540, 12074521, 12611354, 13172055, 13757685, 14369351, 15008212, 15675477, 16372409, 17100326, 17860607, 18654689, 19484076, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396),
(74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 3571900, 3730706, 3896573, 4069815, 4250759, 4439748, 4637139, 4843306, 5058639, 5283546, 5518453, 5763803, 6020062, 6287714, 6567266, 6859246, 7164208, 7482729, 7815411, 8162884, 8525806, 8904863, 9300773, 9714286, 10146183, 10597282, 11068437, 11560540, 12074521, 12611354, 13172055, 13757685, 14369351, 15008212, 15675477, 16372409, 17100326, 17860607, 18654689, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229),
(71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 3571900, 3730706, 3896573, 4069815, 4250759, 4439748, 4637139, 4843306, 5058639, 5283546, 5518453, 5763803, 6020062, 6287714, 6567266, 6859246, 7164208, 7482729, 7815411, 8162884, 8525806, 8904863, 9300773, 9714286, 10146183, 10597282, 11068437, 11560540, 12074521, 12611354, 13172055, 13757685, 14369351, 15008212, 15675477, 16372409, 17100326, 17860607, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197),
(68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 3571900, 3730706, 3896573, 4069815, 4250759, 4439748, 4637139, 4843306, 5058639, 5283546, 5518453, 5763803, 6020062, 6287714, 6567266, 6859246, 7164208, 7482729, 7815411, 8162884, 8525806, 8904863, 9300773, 9714286, 10146183, 10597282, 11068437, 11560540, 12074521, 12611354, 13172055, 13757685, 14369351, 15008212, 15675477, 16372409, 17100326, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295),
(65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 3571900, 3730706, 3896573, 4069815, 4250759, 4439748, 4637139, 4843306, 5058639, 5283546, 5518453, 5763803, 6020062, 6287714, 6567266, 6859246, 7164208, 7482729, 7815411, 8162884, 8525806, 8904863, 9300773, 9714286, 10146183, 10597282, 11068437, 11560540, 12074521, 12611354, 13172055, 13757685, 14369351, 15008212, 15675477, 16372409, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516),
(62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 3571900, 3730706, 3896573, 4069815, 4250759, 4439748, 4637139, 4843306, 5058639, 5283546, 5518453, 5763803, 6020062, 6287714, 6567266, 6859246, 7164208, 7482729, 7815411, 8162884, 8525806, 8904863, 9300773, 9714286, 10146183, 10597282, 11068437, 11560540, 12074521, 12611354, 13172055, 13757685, 14369351, 15008212, 15675477, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855),
(59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 3571900, 3730706, 3896573, 4069815, 4250759, 4439748, 4637139, 4843306, 5058639, 5283546, 5518453, 5763803, 6020062, 6287714, 6567266, 6859246, 7164208, 7482729, 7815411, 8162884, 8525806, 8904863, 9300773, 9714286, 10146183, 10597282, 11068437, 11560540, 12074521, 12611354, 13172055, 13757685, 14369351, 15008212, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307),
(57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 3571900, 3730706, 3896573, 4069815, 4250759, 4439748, 4637139, 4843306, 5058639, 5283546, 5518453, 5763803, 6020062, 6287714, 6567266, 6859246, 7164208, 7482729, 7815411, 8162884, 8525806, 8904863, 9300773, 9714286, 10146183, 10597282, 11068437, 11560540, 12074521, 12611354, 13172055, 13757685, 14369351, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868),
(54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 3571900, 3730706, 3896573, 4069815, 4250759, 4439748, 4637139, 4843306, 5058639, 5283546, 5518453, 5763803, 6020062, 6287714, 6567266, 6859246, 7164208, 7482729, 7815411, 8162884, 8525806, 8904863, 9300773, 9714286, 10146183, 10597282, 11068437, 11560540, 12074521, 12611354, 13172055, 13757685, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533),
(52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 3571900, 3730706, 3896573, 4069815, 4250759, 4439748, 4637139, 4843306, 5058639, 5283546, 5518453, 5763803, 6020062, 6287714, 6567266, 6859246, 7164208, 7482729, 7815411, 8162884, 8525806, 8904863, 9300773, 9714286, 10146183, 10597282, 11068437, 11560540, 12074521, 12611354, 13172055, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297),
(50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 3571900, 3730706, 3896573, 4069815, 4250759, 4439748, 4637139, 4843306, 5058639, 5283546, 5518453, 5763803, 6020062, 6287714, 6567266, 6859246, 7164208, 7482729, 7815411, 8162884, 8525806, 8904863, 9300773, 9714286, 10146183, 10597282, 11068437, 11560540, 12074521, 12611354, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157),
(48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 3571900, 3730706, 3896573, 4069815, 4250759, 4439748, 4637139, 4843306, 5058639, 5283546, 5518453, 5763803, 6020062, 6287714, 6567266, 6859246, 7164208, 7482729, 7815411, 8162884, 8525806, 8904863, 9300773, 9714286, 10146183, 10597282, 11068437, 11560540, 12074521, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107),
(46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 3571900, 3730706, 3896573, 4069815, 4250759, 4439748, 4637139, 4843306, 5058639, 5283546, 5518453, 5763803, 6020062, 6287714, 6567266, 6859246, 7164208, 7482729, 7815411, 8162884, 8525806, 8904863, 9300773, 9714286, 10146183, 10597282, 11068437, 11560540, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145),
(44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 3571900, 3730706, 3896573, 4069815, 4250759, 4439748, 4637139, 4843306, 5058639, 5283546, 5518453, 5763803, 6020062, 6287714, 6567266, 6859246, 7164208, 7482729, 7815411, 8162884, 8525806, 8904863, 9300773, 9714286, 10146183, 10597282, 11068437, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266),
(42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 3571900, 3730706, 3896573, 4069815, 4250759, 4439748, 4637139, 4843306, 5058639, 5283546, 5518453, 5763803, 6020062, 6287714, 6567266, 6859246, 7164208, 7482729, 7815411, 8162884, 8525806, 8904863, 9300773, 9714286, 10146183, 10597282, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468),
(40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 3571900, 3730706, 3896573, 4069815, 4250759, 4439748, 4637139, 4843306, 5058639, 5283546, 5518453, 5763803, 6020062, 6287714, 6567266, 6859246, 7164208, 7482729, 7815411, 8162884, 8525806, 8904863, 9300773, 9714286, 10146183, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746),
(38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 3571900, 3730706, 3896573, 4069815, 4250759, 4439748, 4637139, 4843306, 5058639, 5283546, 5518453, 5763803, 6020062, 6287714, 6567266, 6859246, 7164208, 7482729, 7815411, 8162884, 8525806, 8904863, 9300773, 9714286, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097),
(37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 3571900, 3730706, 3896573, 4069815, 4250759, 4439748, 4637139, 4843306, 5058639, 5283546, 5518453, 5763803, 6020062, 6287714, 6567266, 6859246, 7164208, 7482729, 7815411, 8162884, 8525806, 8904863, 9300773, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518),
(35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 3571900, 3730706, 3896573, 4069815, 4250759, 4439748, 4637139, 4843306, 5058639, 5283546, 5518453, 5763803, 6020062, 6287714, 6567266, 6859246, 7164208, 7482729, 7815411, 8162884, 8525806, 8904863, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007),
(34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 3571900, 3730706, 3896573, 4069815, 4250759, 4439748, 4637139, 4843306, 5058639, 5283546, 5518453, 5763803, 6020062, 6287714, 6567266, 6859246, 7164208, 7482729, 7815411, 8162884, 8525806, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560),
(32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 3571900, 3730706, 3896573, 4069815, 4250759, 4439748, 4637139, 4843306, 5058639, 5283546, 5518453, 5763803, 6020062, 6287714, 6567266, 6859246, 7164208, 7482729, 7815411, 8162884, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175),
(31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 3571900, 3730706, 3896573, 4069815, 4250759, 4439748, 4637139, 4843306, 5058639, 5283546, 5518453, 5763803, 6020062, 6287714, 6567266, 6859246, 7164208, 7482729, 7815411, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848),
(29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 3571900, 3730706, 3896573, 4069815, 4250759, 4439748, 4637139, 4843306, 5058639, 5283546, 5518453, 5763803, 6020062, 6287714, 6567266, 6859246, 7164208, 7482729, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579),
(28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 3571900, 3730706, 3896573, 4069815, 4250759, 4439748, 4637139, 4843306, 5058639, 5283546, 5518453, 5763803, 6020062, 6287714, 6567266, 6859246, 7164208, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363),
(27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 3571900, 3730706, 3896573, 4069815, 4250759, 4439748, 4637139, 4843306, 5058639, 5283546, 5518453, 5763803, 6020062, 6287714, 6567266, 6859246, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199),
(26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 3571900, 3730706, 3896573, 4069815, 4250759, 4439748, 4637139, 4843306, 5058639, 5283546, 5518453, 5763803, 6020062, 6287714, 6567266, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085),
(25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 3571900, 3730706, 3896573, 4069815, 4250759, 4439748, 4637139, 4843306, 5058639, 5283546, 5518453, 5763803, 6020062, 6287714, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018),
(24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 3571900, 3730706, 3896573, 4069815, 4250759, 4439748, 4637139, 4843306, 5058639, 5283546, 5518453, 5763803, 6020062, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996),
(22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 3571900, 3730706, 3896573, 4069815, 4250759, 4439748, 4637139, 4843306, 5058639, 5283546, 5518453, 5763803, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018),
(22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 3571900, 3730706, 3896573, 4069815, 4250759, 4439748, 4637139, 4843306, 5058639, 5283546, 5518453, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082),
(21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 3571900, 3730706, 3896573, 4069815, 4250759, 4439748, 4637139, 4843306, 5058639, 5283546, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186),
(20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 3571900, 3730706, 3896573, 4069815, 4250759, 4439748, 4637139, 4843306, 5058639, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327),
(19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 3571900, 3730706, 3896573, 4069815, 4250759, 4439748, 4637139, 4843306, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506),
(18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 3571900, 3730706, 3896573, 4069815, 4250759, 4439748, 4637139, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719),
(17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 3571900, 3730706, 3896573, 4069815, 4250759, 4439748, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966),
(16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 3571900, 3730706, 3896573, 4069815, 4250759, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245),
(16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 3571900, 3730706, 3896573, 4069815, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555),
(15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 3571900, 3730706, 3896573, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894),
(14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 3571900, 3730706, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262),
(14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 3571900, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656),
(13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 3419853, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077),
(13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 3274279, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522),
(12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 3134901, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990),
(11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 3001456, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482),
(11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 2873692, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995),
(10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 2751366, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529),
(10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 2634248, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083),
(10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 2522114, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656),
(9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 2414754, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247),
(9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 2311964, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856),
(8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 2213550, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481),
(8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 2119325, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123),
(8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 2029111, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780),
(7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 1942737, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451),
(7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 1860039, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137),
(7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 1780862, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836),
(6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 1705055, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548),
(6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 1632476, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273),
(6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 1562985, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010),
(6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 1496453, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757),
(5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 1432753, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516),
(5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 1371764, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285),
(5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 1313372, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064),
(5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 1257465, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853),
(4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 1203938, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651),
(4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 1152689, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458),
(4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 1103622, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273),
(4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 1056644, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096),
(4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 1011665, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927),
(3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 968601, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766),
(3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 927370, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611),
(3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 887895, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464),
(3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 850099, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323),
(3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 813913, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188),
(3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 779267, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059),
(3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 746095, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936),
(2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 714336, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819),
(2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 683928, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707),
(2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 654815, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600),
(2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 626942, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498),
(2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 600254, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401),
(2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 574703, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308),
(2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 550240, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220),
(2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 526817, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136),
(2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 504392, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056),
(2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 482921, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979),
(1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 462365, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907),
(1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 442683, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838),
(1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 423839, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773),
(1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 405798, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711),
(1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 388524, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652),
(1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 371985, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596),
(1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 356151, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544),
(1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 340991, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494),
(1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 326476, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447),
(1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 312578, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403),
(1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 299273, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361),
(1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 286534, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323),
(1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 274337, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286),
(1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 262659, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252),
(1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 251478, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221),
(1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 240774, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191),
(1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 230525, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164),
(1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 220712, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139),
(1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 211317, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117),
(1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 202322, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096),
(1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 193709, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078),
(1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 185464, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061),
(1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 177569, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034, 1047),
(1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 170011, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024, 1034),
(1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 162774, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015, 1024),
(1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 155845, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009, 1015),
(1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 149211, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004, 1009),
(1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 142860, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001, 1004),
(1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 136779, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000, 1001),
(1001, 1004, 1009, 1015, 1024, 1034, 1047, 1061, 1078, 1096, 1117, 1139, 1164, 1191, 1221, 1252, 1286, 1323, 1361, 1403, 1447, 1494, 1544, 1596, 1652, 1711, 1773, 1838, 1907, 1979, 2056, 2136, 2220, 2308, 2401, 2498, 2600, 2707, 2819, 2936, 3059, 3188, 3323, 3464, 3611, 3766, 3927, 4096, 4273, 4458, 4651, 4853, 5064, 5285, 5516, 5757, 6010, 6273, 6548, 6836, 7137, 7451, 7780, 8123, 8481, 8856, 9247, 9656, 10083, 10529, 10995, 11482, 11990, 12522, 13077, 13656, 14262, 14894, 15555, 16245, 16966, 17719, 18506, 19327, 20186, 21082, 22018, 22996, 24018, 25085, 26199, 27363, 28579, 29848, 31175, 32560, 34007, 35518, 37097, 38746, 40468, 42266, 44145, 46107, 48157, 50297, 52533, 54868, 57307, 59855, 62516, 65295, 68197, 71229, 74396, 77703, 81157, 84765, 88534, 92470, 96581, 100875, 105359, 110043, 114936, 120045, 125382, 130957, 125382, 120045, 114936, 110043, 105359, 100875, 96581, 92470, 88534, 84765, 81157, 77703, 74396, 71229, 68197, 65295, 62516, 59855, 57307, 54868, 52533, 50297, 48157, 46107, 44145, 42266, 40468, 38746, 37097, 35518, 34007, 32560, 31175, 29848, 28579, 27363, 26199, 25085, 24018, 22996, 22018, 21082, 20186, 19327, 18506, 17719, 16966, 16245, 15555, 14894, 14262, 13656, 13077, 12522, 11990, 11482, 10995, 10529, 10083, 9656, 9247, 8856, 8481, 8123, 7780, 7451, 7137, 6836, 6548, 6273, 6010, 5757, 5516, 5285, 5064, 4853, 4651, 4458, 4273, 4096, 3927, 3766, 3611, 3464, 3323, 3188, 3059, 2936, 2819, 2707, 2600, 2498, 2401, 2308, 2220, 2136, 2056, 1979, 1907, 1838, 1773, 1711, 1652, 1596, 1544, 1494, 1447, 1403, 1361, 1323, 1286, 1252, 1221, 1191, 1164, 1139, 1117, 1096, 1078, 1061, 1047, 1034, 1024, 1015, 1009, 1004, 1001, 1000)

);

type calo_calo_cos_dphi_lut_array is array (0 to 143, 0 to 143) of integer;
constant CALO_CALO_COS_DPHI_LUT: calo_calo_cos_dphi_lut_array := (

(1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999),
(999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996),
(996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991),
(991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985),
(985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976),
(976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966),
(966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954),
(954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940),
(940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924),
(924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906),
(906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887),
(887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866),
(866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843),
(843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819),
(819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793),
(793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766),
(766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737),
(737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707),
(707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676),
(676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643),
(643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609),
(609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574),
(574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537),
(537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500),
(500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462),
(462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423),
(423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383),
(383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342),
(342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301),
(301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259),
(259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216),
(216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174),
(174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131),
(131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87),
(87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44),
(44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0),
(0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44),
(-44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87),
(-87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131),
(-131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174),
(-174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216),
(-216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259),
(-259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301),
(-301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342),
(-342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383),
(-383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423),
(-423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462),
(-462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500),
(-500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537),
(-537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574),
(-574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609),
(-609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643),
(-643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676),
(-676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707),
(-707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737),
(-737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766),
(-766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793),
(-793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819),
(-819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843),
(-843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866),
(-866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887),
(-887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906),
(-906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924),
(-924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940),
(-940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954),
(-954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966),
(-966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976),
(-976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985),
(-985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991),
(-991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996),
(-996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999),
(-999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000),
(-1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999),
(-999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996),
(-996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991),
(-991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985),
(-985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976),
(-976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966),
(-966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954),
(-954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940),
(-940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924),
(-924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906),
(-906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887),
(-887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866),
(-866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843),
(-843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819),
(-819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793),
(-793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766),
(-766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737),
(-737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707),
(-707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676),
(-676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643),
(-643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609),
(-609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574),
(-574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537),
(-537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500),
(-500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462),
(-462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423),
(-423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383),
(-383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342),
(-342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301),
(-301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259),
(-259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216),
(-216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174),
(-174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131),
(-131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87),
(-87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44),
(-44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0),
(0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44),
(44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87),
(87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131),
(131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174),
(174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216),
(216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259),
(259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301),
(301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342),
(342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383),
(383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423),
(423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462),
(462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500),
(500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537),
(537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574),
(574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609),
(609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643),
(643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676),
(676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707),
(707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737),
(737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766),
(766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793),
(793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819),
(819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843),
(843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866),
(866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887),
(887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924, 906),
(906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940, 924),
(924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954, 940),
(940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966, 954),
(954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976, 966),
(966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985, 976),
(976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991, 985),
(985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996, 991),
(991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999, 996),
(996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000, 999),
(999, 996, 991, 985, 976, 966, 954, 940, 924, 906, 887, 866, 843, 819, 793, 766, 737, 707, 676, 643, 609, 574, 537, 500, 462, 423, 383, 342, 301, 259, 216, 174, 131, 87, 44, 0, -44, -87, -131, -174, -216, -259, -301, -342, -383, -423, -462, -500, -537, -574, -609, -643, -676, -707, -737, -766, -793, -819, -843, -866, -887, -906, -924, -940, -954, -966, -976, -985, -991, -996, -999, -1000, -999, -996, -991, -985, -976, -966, -954, -940, -924, -906, -887, -866, -843, -819, -793, -766, -737, -707, -676, -643, -609, -574, -537, -500, -462, -423, -383, -342, -301, -259, -216, -174, -131, -87, -44, 0, 44, 87, 131, 174, 216, 259, 301, 342, 383, 423, 462, 500, 537, 574, 609, 643, 676, 707, 737, 766, 793, 819, 843, 866, 887, 906, 924, 940, 954, 966, 976, 985, 991, 996, 999, 1000)

);

end package;
