
library ieee;
use ieee.std_logic_1164.all;

package algo_pre_scaler_fractional_tb_pkg is

    constant PRESCALE_FACTOR_VAL : std_logic_vector(31 downto 0) := X"13000001"; -- actual factor for test = 1.95

end algo_pre_scaler_fractional_tb_pkg;
