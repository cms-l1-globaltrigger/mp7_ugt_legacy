-- Description:
-- Package for deltaR LUT for invariant mass divided by deltaR. 
-- Calculation of values: 1/DR**2 rounded with precision 5 and multiplicated with 10**5.
-- These values are used for formular: invariant mass * 1/DR**2

-- Version history:
-- HB 2020-04-22: first design

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

use work.gtl_pkg.all;

package delta_r_lut_pkg is

constant CALO_DETA_BINS : positive := 230;
constant CALO_DPHI_BINS : positive := 144;

constant MAX_WIDTH_MASS_DIV_DR_LIMIT_VECTOR : positive := 80;

constant CALO_INV_DR_SQ_LUT_MAX_VAL : natural := 52847140;
constant CALO_INV_DR_SQ_VECTOR_WIDTH : natural := 26; -- => log2(CALO_INV_DR_SQ_LUT_MAX_VAL)
constant EG_EG_INV_DR_SQ_VECTOR_WIDTH : natural := CALO_INV_DR_SQ_VECTOR_WIDTH;
constant EG_JET_INV_DR_SQ_VECTOR_WIDTH : natural := CALO_INV_DR_SQ_VECTOR_WIDTH;
constant EG_TAU_INV_DR_SQ_VECTOR_WIDTH : natural := CALO_INV_DR_SQ_VECTOR_WIDTH;
constant JET_JET_INV_DR_SQ_VECTOR_WIDTH : natural := CALO_INV_DR_SQ_VECTOR_WIDTH;
constant JET_TAU_INV_DR_SQ_VECTOR_WIDTH : natural := CALO_INV_DR_SQ_VECTOR_WIDTH;
constant TAU_TAU_INV_DR_SQ_VECTOR_WIDTH : natural := CALO_INV_DR_SQ_VECTOR_WIDTH;

type calo_inv_dr_sq_vector_array is array (natural range <>, natural range <>) of std_logic_vector(CALO_INV_DR_SQ_VECTOR_WIDTH-1 downto 0);

-- Value of first LUT address has to be defined, it's the division by 0 (actually = 0) !!! 

type calo_inv_dr_sq_lut_array is array (0 to CALO_DETA_BINS-1, 0 to CALO_DPHI_BINS-1) of natural range 0 to CALO_INV_DR_SQ_LUT_MAX_VAL;
constant CALO_INV_DR_SQ_LUT : calo_inv_dr_sq_lut_array := (
(0, 52524902, 13131225, 5836100, 3282806, 2100996, 1459025, 1071937, 820702, 648456, 525249, 434090, 364756, 310798, 267984, 233443,
205175, 181747, 162114, 145498, 131312, 119104, 108522, 99291, 91189, 84040, 77700, 72051, 66996, 62455, 58360, 54657,
51293, 48232, 45437, 42877, 40528, 38367, 36375, 34533, 32828, 31246, 29776, 28407, 27131, 25938, 24823, 23778,
22797, 21876, 21010, 20194, 19425, 18699, 18013, 17364, 16749, 16166, 15614, 15089, 14590, 14116, 13664, 13234,
12823, 12432, 12058, 11701, 11359, 11032, 10719, 10420, 10132, 9856, 9592, 9338, 9094, 8859, 8633, 8416,
8207, 8006, 7811, 7624, 7444, 7270, 7102, 6938, 6783, 6630, 6485, 6343, 6206, 6073, 5944, 5820,
5699, 5582, 5469, 5359, 5252, 5149, 5049, 4951, 4856, 4764, 4675, 4588, 4503, 4421, 4341, 4263,
4187, 4113, 4041, 3972, 3903, 3837, 3771, 3709, 3648, 3588, 3529, 3472, 3416, 3361, 3308, 3257,
3206, 3156, 3108, 3061, 3015, 2969, 2925, 2882, 2840, 2798, 2758, 2719, 2680, 2642, 2605, 2569),
(52847140, 26342764, 10517807, 5255695, 3090809, 2020662, 1419826, 1050626, 808151, 640595, 520080, 430553, 362256, 308981, 266632, 232417,
204382, 181124, 161618, 145099, 130987, 118836, 108300, 99105, 91032, 83906, 77585, 71953, 66911, 62382, 58297, 54600,
51244, 48188, 45398, 42843, 40497, 38340, 36350, 34511, 32808, 31228, 29759, 28392, 27117, 25924, 24811, 23767,
22787, 21867, 21002, 20186, 19418, 18692, 18007, 17358, 16744, 16162, 15609, 15085, 14585, 14112, 13661, 13230,
12820, 12429, 12055, 11698, 11357, 11030, 10717, 10417, 10130, 9855, 9590, 9336, 9092, 8857, 8632, 8415,
8206, 8004, 7810, 7623, 7443, 7269, 7101, 6938, 6782, 6630, 6483, 6342, 6205, 6072, 5944, 5819,
5699, 5582, 5468, 5359, 5252, 5148, 5048, 4951, 4856, 4764, 4674, 4587, 4503, 4421, 4341, 4263,
4187, 4113, 4041, 3971, 3903, 3837, 3771, 3709, 3647, 3587, 3529, 3472, 3416, 3361, 3308, 3256,
3206, 3156, 3108, 3061, 3014, 2969, 2925, 2882, 2840, 2798, 2758, 2718, 2680, 2642, 2605, 2568),
(13211785, 10556475, 6585691, 4047972, 2629452, 1812728, 1313924, 991492, 772702, 618117, 505166, 420281, 354956, 303655, 262657, 229391,
202037, 179281, 160149, 143913, 130020, 118039, 107637, 98550, 90564, 83509, 77245, 71660, 66658, 62161, 58104, 54430,
51095, 48057, 45281, 42739, 40405, 38256, 36275, 34443, 32747, 31172, 29709, 28346, 27075, 25887, 24776, 23735,
22758, 21840, 20977, 20163, 19396, 18672, 17988, 17341, 16728, 16147, 15595, 15072, 14574, 14101, 13650, 13221,
12811, 12420, 12047, 11690, 11349, 11023, 10711, 10411, 10124, 9849, 9585, 9331, 9087, 8853, 8628, 8411,
8202, 8001, 7807, 7620, 7439, 7266, 7098, 6936, 6779, 6628, 6481, 6340, 6203, 6070, 5942, 5817,
5697, 5580, 5467, 5357, 5250, 5147, 5047, 4949, 4854, 4762, 4673, 4586, 4502, 4419, 4339, 4262,
4186, 4112, 4040, 3970, 3902, 3836, 3771, 3708, 3647, 3587, 3528, 3471, 3415, 3361, 3308, 3256,
3205, 3156, 3107, 3060, 3014, 2969, 2925, 2881, 2839, 2798, 2758, 2718, 2679, 2641, 2604, 2568),
(5871904, 5281474, 4057504, 2926974, 2105618, 1547348, 1168645, 906459, 720061, 583966, 482123, 404208, 343423, 295175, 256287, 224518,
198248, 176291, 157758, 141980, 128440, 116736, 106553, 97640, 89795, 82854, 76685, 71177, 66240, 61798, 57787, 54152,
50849, 47839, 45088, 42567, 40251, 38118, 36151, 34331, 32645, 31080, 29626, 28270, 27006, 25824, 24718, 23682,
22709, 21795, 20935, 20125, 19361, 18639, 17958, 17312, 16701, 16122, 15572, 15050, 14554, 14082, 13632, 13203,
12795, 12406, 12033, 11678, 11337, 11012, 10700, 10401, 10115, 9840, 9576, 9323, 9080, 8846, 8621, 8404,
8196, 7994, 7801, 7615, 7435, 7260, 7093, 6931, 6775, 6623, 6476, 6336, 6199, 6067, 5938, 5814,
5694, 5577, 5464, 5354, 5248, 5144, 5044, 4947, 4852, 4760, 4671, 4584, 4500, 4418, 4338, 4260,
4184, 4111, 4039, 3969, 3901, 3835, 3769, 3707, 3645, 3585, 3527, 3470, 3413, 3360, 3307, 3255,
3204, 3155, 3106, 3059, 3013, 2968, 2924, 2881, 2838, 2797, 2757, 2717, 2679, 2641, 2604, 2567),
(3302946, 3107534, 2639119, 2109227, 1646423, 1284151, 1011993, 809290, 657363, 542039, 453182, 383667, 328481, 284068, 247873, 218034,
193176, 172268, 154529, 139359, 126291, 114958, 105070, 96393, 88739, 81955, 75914, 70512, 65664, 61295, 57348, 53767,
50509, 47538, 44820, 42328, 40037, 37927, 35978, 34176, 32505, 30953, 29509, 28165, 26910, 25735, 24638, 23608,
22641, 21732, 20877, 20071, 19311, 18594, 17915, 17273, 16665, 16088, 15540, 15020, 14526, 14055, 13608, 13181,
12774, 12385, 12014, 11659, 11320, 10996, 10685, 10387, 10101, 9827, 9564, 9311, 9069, 8835, 8611, 8395,
8187, 7986, 7793, 7607, 7427, 7253, 7087, 6925, 6769, 6618, 6472, 6331, 6194, 6062, 5934, 5810,
5689, 5573, 5460, 5350, 5244, 5141, 5041, 4944, 4849, 4757, 4668, 4581, 4497, 4415, 4335, 4258,
4182, 4108, 4037, 3966, 3898, 3833, 3768, 3705, 3644, 3583, 3524, 3468, 3413, 3358, 3305, 3253,
3203, 3153, 3105, 3058, 3012, 2967, 2923, 2880, 2837, 2796, 2756, 2716, 2678, 2640, 2603, 2567),
(2113886, 2032103, 1820774, 1551808, 1285876, 1053711, 863221, 711261, 591180, 496232, 420712, 360136, 311079, 270960, 237833, 210228,
187023, 167358, 150567, 136129, 123632, 112751, 103223, 94836, 87418, 80826, 74945, 69676, 64937, 60663, 56793, 53279,
50078, 47156, 44481, 42025, 39766, 37683, 35759, 33978, 32326, 30791, 29362, 28031, 26787, 25624, 24535, 23513,
22554, 21652, 20803, 20003, 19248, 18535, 17860, 17222, 16617, 16044, 15498, 14982, 14490, 14022, 13576, 13150,
12745, 12359, 11990, 11636, 11298, 10975, 10665, 10368, 10084, 9811, 9549, 9297, 9055, 8822, 8598, 8383,
8175, 7975, 7783, 7597, 7418, 7245, 7078, 6916, 6761, 6610, 6465, 6324, 6188, 6056, 5928, 5804,
5684, 5568, 5455, 5346, 5239, 5136, 5037, 4939, 4845, 4753, 4664, 4578, 4494, 4412, 4332, 4254,
4179, 4105, 4034, 3964, 3896, 3830, 3766, 3703, 3641, 3581, 3522, 3466, 3411, 3356, 3302, 3252,
3200, 3152, 3103, 3056, 3010, 2965, 2921, 2878, 2836, 2795, 2754, 2715, 2676, 2639, 2602, 2565),
(1467976, 1428064, 1320368, 1172942, 1014376, 864174, 731743, 619540, 526405, 449775, 386837, 335022, 292161, 256494, 226615, 201413,
180015, 161724, 145992, 132378, 120531, 110166, 101052, 93001, 85856, 79489, 73794, 68680, 64071, 59907, 56130, 52695,
49562, 46698, 44073, 41661, 39440, 37390, 35495, 33739, 32110, 30595, 29184, 27868, 26638, 25488, 24410, 23399,
22449, 21555, 20714, 19920, 19171, 18464, 17794, 17161, 16560, 15989, 15448, 14936, 14446, 13980, 13538, 13116,
12712, 12328, 11960, 11608, 11272, 10950, 10642, 10346, 10063, 9791, 9530, 9279, 9038, 8806, 8583, 8368,
8161, 7962, 7770, 7585, 7406, 7234, 7068, 6907, 6751, 6601, 6456, 6315, 6180, 6048, 5920, 5797,
5677, 5561, 5449, 5340, 5234, 5131, 5031, 4934, 4840, 4749, 4660, 4573, 4489, 4408, 4328, 4251,
4175, 4102, 4031, 3961, 3893, 3827, 3762, 3700, 3639, 3579, 3520, 3463, 3408, 3354, 3300, 3249,
3198, 3150, 3101, 3054, 3008, 2963, 2919, 2876, 2834, 2793, 2753, 2714, 2675, 2637, 2600, 2564),
(1078513, 1056813, 996654, 910291, 811807, 712673, 620120, 537607, 466054, 404968, 353224, 309514, 272572, 241271, 214649, 191906,
172382, 155537, 140930, 128203, 117060, 107259, 98601, 90921, 84080, 77965, 72478, 67539, 63078, 59036, 55365, 52020,
48965, 46168, 43600, 41238, 39061, 37049, 35188, 33462, 31857, 30366, 28976, 27678, 26465, 25329, 24264, 23265,
22325, 21441, 20608, 19823, 19081, 18380, 17717, 17088, 16493, 15928, 15391, 14881, 14396, 13933, 13493, 13073,
12673, 12290, 11925, 11575, 11241, 10921, 10614, 10320, 10038, 9767, 9507, 9258, 9018, 8787, 8565, 8351,
8144, 7947, 7754, 7571, 7393, 7221, 7055, 6895, 6740, 6591, 6446, 6306, 6170, 6039, 5912, 5789,
5669, 5554, 5441, 5333, 5227, 5125, 5025, 4928, 4834, 4743, 4655, 4568, 4484, 4403, 4323, 4246,
4171, 4098, 4027, 3957, 3889, 3823, 3759, 3696, 3635, 3576, 3517, 3461, 3404, 3351, 3298, 3247,
3196, 3147, 3099, 3052, 3006, 2961, 2917, 2874, 2832, 2791, 2751, 2712, 2673, 2636, 2599, 2562),
(825737, 812956, 776883, 723386, 659780, 592767, 527307, 466432, 411606, 363218, 321038, 284519, 252998, 225807, 202323, 181993,
164341, 148960, 135510, 123702, 113296, 104090, 95917, 88633, 82120, 76277, 71017, 66268, 61968, 58064, 54508, 51263,
48294, 45570, 43067, 40761, 38632, 36664, 34840, 33147, 31573, 30107, 28740, 27461, 26268, 25147, 24098, 23112,
22185, 21312, 20489, 19712, 18978, 18285, 17628, 17006, 16416, 15856, 15323, 14818, 14337, 13879, 13442, 13025,
12627, 12248, 11885, 11537, 11205, 10887, 10582, 10290, 10009, 9740, 9482, 9233, 8995, 8765, 8544, 8331,
8126, 7929, 7738, 7555, 7377, 7206, 7041, 6882, 6727, 6578, 6433, 6294, 6159, 6029, 5902, 5779,
5660, 5545, 5433, 5325, 5219, 5117, 5018, 4921, 4828, 4737, 4648, 4562, 4479, 4397, 4318, 4241,
4166, 4093, 4022, 3953, 3885, 3819, 3755, 3692, 3632, 3572, 3513, 3456, 3402, 3348, 3295, 3243,
3193, 3144, 3096, 3049, 3004, 2959, 2915, 2872, 2830, 2789, 2749, 2710, 2671, 2634, 2597, 2561),
(652434, 644429, 621552, 586830, 544265, 497837, 450833, 405579, 363479, 325219, 290987, 260662, 233958, 210516, 189959, 171928,
156089, 142149, 129848, 118968, 109312, 100718, 93046, 86176, 80007, 74450, 69431, 64885, 60757, 56999, 53569, 50432,
47555, 44912, 42478, 40233, 38158, 36236, 34454, 32797, 31255, 29818, 28476, 27222, 26046, 24946, 23913, 22942,
22028, 21167, 20354, 19588, 18863, 18178, 17529, 16913, 16330, 15776, 15248, 14748, 14271, 13816, 13383, 12971,
12576, 12199, 11839, 11495, 11165, 10849, 10546, 10256, 9977, 9710, 9453, 9206, 8969, 8740, 8521, 8309,
8105, 7908, 7718, 7536, 7360, 7190, 7025, 6866, 6712, 6564, 6421, 6282, 6147, 6017, 5891, 5768,
5650, 5535, 5424, 5315, 5211, 5109, 5010, 4914, 4820, 4730, 4641, 4556, 4472, 4391, 4312, 4235,
4161, 4088, 4016, 3948, 3880, 3815, 3751, 3688, 3626, 3568, 3510, 3453, 3398, 3343, 3292, 3240,
3190, 3141, 3093, 3046, 3001, 2956, 2912, 2869, 2827, 2787, 2746, 2707, 2669, 2631, 2595, 2559),
(528471, 523207, 508026, 484591, 455194, 422259, 387952, 353965, 321469, 291174, 263428, 238327, 215804, 195703, 177815, 161919,
147795, 135237, 124058, 114087, 105178, 97198, 90034, 83586, 77770, 72509, 67740, 63405, 59458, 55854, 52557, 49534,
46756, 44198, 41840, 39660, 37642, 35770, 34032, 32415, 30908, 29502, 28188, 26958, 25806, 24725, 23709, 22754,
21855, 21007, 20207, 19451, 18736, 18060, 17419, 16811, 16234, 15687, 15165, 14670, 14198, 13749, 13320, 12910,
12520, 12146, 11789, 11447, 11120, 10807, 10506, 10218, 9942, 9676, 9421, 9176, 8940, 8713, 8495, 8284,
8082, 7886, 7698, 7516, 7341, 7171, 7008, 6850, 6697, 6549, 6406, 6268, 6134, 6004, 5878, 5757,
5639, 5524, 5413, 5305, 5201, 5099, 5001, 4905, 4812, 4722, 4634, 4548, 4465, 4384, 4306, 4229,
4154, 4082, 4011, 3941, 3875, 3809, 3746, 3683, 3623, 3563, 3506, 3449, 3394, 3340, 3288, 3237,
3187, 3138, 3090, 3043, 2997, 2953, 2909, 2866, 2825, 2784, 2744, 2705, 2666, 2629, 2592, 2556),
(436753, 433151, 422694, 406344, 385469, 361587, 336133, 310317, 285055, 260977, 238465, 217709, 198761, 181582, 166080, 152130,
139597, 128340, 118229, 109139, 100959, 93584, 86924, 80899, 75438, 70478, 65964, 61848, 58086, 54642, 51482, 48577,
45903, 43435, 41155, 39044, 37087, 35269, 33578, 32002, 30533, 29160, 27876, 26672, 25544, 24484, 23488, 22550,
21666, 20833, 20046, 19302, 18598, 17931, 17299, 16700, 16130, 15589, 15075, 14585, 14119, 13674, 13250, 12845,
12458, 12088, 11734, 11396, 11071, 10761, 10463, 10177, 9902, 9639, 9386, 9142, 8908, 8683, 8466, 8257,
8056, 7861, 7674, 7494, 7319, 7151, 6988, 6831, 6679, 6532, 6390, 6252, 6119, 5990, 5865, 5743,
5626, 5512, 5401, 5294, 5190, 5089, 4991, 4895, 4803, 4713, 4625, 4540, 4457, 4377, 4298, 4222,
4147, 4075, 4005, 3936, 3869, 3803, 3740, 3678, 3617, 3558, 3501, 3444, 3390, 3336, 3284, 3232,
3182, 3134, 3086, 3039, 2994, 2949, 2906, 2863, 2821, 2781, 2741, 2702, 2663, 2626, 2589, 2554),
(366994, 364448, 357016, 345282, 330092, 312421, 293235, 273394, 253594, 234358, 216042, 198866, 182936, 168283, 154885, 142683,
131601, 121551, 112444, 104190, 96709, 89921, 83755, 78148, 73040, 68381, 64123, 60227, 56654, 53372, 50354, 47572,
45004, 42630, 40431, 38392, 36498, 34736, 33094, 31563, 30133, 28795, 27541, 26366, 25263, 24226, 23250, 22331,
21464, 20646, 19872, 19141, 18448, 17792, 17170, 16579, 16017, 15484, 14976, 14493, 14032, 13593, 13174, 12773,
12391, 12025, 11674, 11339, 11018, 10710, 10415, 10132, 9860, 9599, 9348, 9106, 8874, 8650, 8435, 8227,
8026, 7835, 7649, 7469, 7296, 7129, 6967, 6811, 6660, 6512, 6372, 6235, 6102, 5974, 5850, 5729,
5612, 5499, 5389, 5282, 5178, 5078, 4980, 4885, 4793, 4703, 4616, 4531, 4449, 4368, 4290, 4214,
4140, 4068, 3998, 3929, 3862, 3796, 3734, 3672, 3612, 3553, 3495, 3438, 3385, 3331, 3279, 3228,
3178, 3129, 3082, 3035, 2990, 2946, 2902, 2860, 2818, 2777, 2738, 2699, 2660, 2623, 2587, 2551),
(312705, 310854, 305431, 296802, 285509, 272193, 257513, 242084, 226430, 210969, 196011, 181766, 168365, 155874, 144311, 133662,
123888, 114942, 106765, 99297, 92478, 86252, 80563, 75362, 70601, 66238, 62236, 58558, 55174, 52058, 49182, 46525,
44066, 41787, 39672, 37707, 35878, 34174, 32584, 31099, 29709, 28408, 27187, 26040, 24965, 23951, 22997, 22097,
21248, 20446, 19687, 18969, 18289, 17644, 17032, 16450, 15898, 15372, 14871, 14394, 13940, 13506, 13092, 12695,
12318, 11957, 11610, 11279, 10961, 10656, 10364, 10084, 9814, 9555, 9306, 9067, 8837, 8615, 8401, 8196,
7997, 7806, 7621, 7443, 7271, 7105, 6944, 6789, 6639, 6493, 6353, 6217, 6085, 5957, 5834, 5714,
5597, 5485, 5375, 5269, 5166, 5066, 4968, 4874, 4782, 4693, 4606, 4521, 4439, 4359, 4281, 4206,
4132, 4059, 3990, 3922, 3855, 3791, 3726, 3666, 3606, 3547, 3490, 3434, 3379, 3326, 3274, 3223,
3173, 3125, 3077, 3031, 2986, 2941, 2898, 2856, 2814, 2774, 2734, 2695, 2657, 2620, 2583, 2548),
(269628, 268251, 264203, 257722, 249164, 238960, 227572, 215438, 202952, 190442, 178168, 166321, 155030, 144377, 134402, 125116,
116514, 108566, 101242, 94502, 88306, 82612, 77378, 72568, 68143, 64070, 60318, 56857, 53662, 50709, 47976, 45444,
43095, 40913, 38884, 36994, 35233, 33588, 32051, 30612, 29265, 28000, 26815, 25700, 24650, 23662, 22730, 21851,
21020, 20235, 19491, 18787, 18120, 17486, 16885, 16313, 15769, 15251, 14759, 14288, 13841, 13414, 13005, 12615,
12241, 11884, 11542, 11214, 10900, 10599, 10310, 10032, 9765, 9509, 9262, 9025, 8797, 8577, 8365, 8161,
7965, 7775, 7592, 7414, 7244, 7079, 6920, 6765, 6616, 6472, 6332, 6197, 6066, 5939, 5816, 5697,
5581, 5469, 5360, 5255, 5152, 5053, 4956, 4862, 4770, 4681, 4595, 4511, 4429, 4350, 4272, 4197,
4123, 4052, 3982, 3914, 3848, 3783, 3719, 3658, 3599, 3540, 3483, 3428, 3373, 3320, 3268, 3218,
3168, 3120, 3073, 3026, 2981, 2937, 2894, 2852, 2810, 2770, 2730, 2691, 2653, 2616, 2580, 2544),
(234876, 233831, 230749, 225789, 219193, 211259, 202308, 192661, 182614, 172423, 162300, 152410, 142875, 133778, 125170, 117079,
109512, 102462, 95913, 89843, 84225, 79029, 74227, 69789, 65687, 61894, 58385, 55137, 52127, 49336, 46746, 44339,
42100, 40015, 38072, 36258, 34564, 32980, 31497, 30107, 28802, 27578, 26426, 25341, 24321, 23359, 22450, 21592,
20780, 20012, 19285, 18595, 17941, 17320, 16730, 16167, 15634, 15125, 14641, 14177, 13737, 13316, 12913, 12528,
12160, 11807, 11469, 11146, 10835, 10537, 10252, 9977, 9713, 9459, 9215, 8981, 8755, 8537, 8327, 8125,
7930, 7742, 7560, 7385, 7215, 7052, 6893, 6740, 6592, 6449, 6310, 6176, 6046, 5920, 5798, 5679,
5564, 5453, 5345, 5240, 5138, 5039, 4942, 4849, 4758, 4669, 4583, 4500, 4418, 4339, 4262, 4187,
4114, 4043, 3973, 3905, 3839, 3775, 3713, 3651, 3592, 3534, 3477, 3420, 3367, 3314, 3262, 3212,
3163, 3115, 3067, 3021, 2976, 2932, 2889, 2847, 2806, 2766, 2726, 2687, 2650, 2613, 2576, 2541),
(206434, 205626, 203239, 199382, 194221, 187966, 180847, 173099, 164945, 156586, 148192, 139903, 131827, 124044, 116608, 109555,
102901, 96653, 90805, 85345, 80259, 75528, 71130, 67044, 63249, 59724, 56452, 53408, 50581, 47949, 45498, 43215,
41085, 39097, 37240, 35503, 33877, 32354, 30925, 29584, 28324, 27138, 26023, 24971, 23979, 23043, 22158, 21322,
20530, 19780, 19069, 18395, 17754, 17146, 16567, 16016, 15492, 14992, 14516, 14061, 13627, 13211, 12816, 12437,
12073, 11726, 11393, 11073, 10767, 10473, 10190, 9919, 9658, 9407, 9166, 8934, 8710, 8494, 8287, 8086,
7893, 7707, 7527, 7353, 7185, 7023, 6866, 6714, 6567, 6425, 6286, 6154, 6025, 5899, 5778, 5660,
5546, 5435, 5328, 5224, 5122, 5024, 4928, 4835, 4745, 4657, 4571, 4488, 4407, 4328, 4252, 4177,
4104, 4033, 3964, 3896, 3830, 3767, 3705, 3644, 3583, 3526, 3470, 3413, 3360, 3308, 3256, 3206,
3157, 3109, 3062, 3016, 2971, 2927, 2884, 2842, 2801, 2761, 2722, 2683, 2645, 2609, 2572, 2537),
(182862, 182228, 180351, 177307, 173214, 168221, 162496, 156214, 149542, 142639, 135640, 128663, 121800, 115126, 108694, 102540,
96689, 91151, 85932, 81027, 76429, 72126, 68105, 64349, 60846, 57577, 54530, 51686, 49032, 46555, 44241, 42079,
40057, 38166, 36394, 34733, 33176, 31713, 30340, 29048, 27832, 26686, 25606, 24588, 23625, 22716, 21856, 21042,
20270, 19539, 18845, 18186, 17560, 16964, 16397, 15858, 15344, 14853, 14385, 13938, 13511, 13103, 12714, 12341,
11983, 11641, 11312, 10997, 10695, 10405, 10126, 9858, 9600, 9352, 9114, 8884, 8663, 8450, 8244, 8046,
7854, 7670, 7492, 7319, 7153, 6992, 6836, 6686, 6540, 6399, 6261, 6130, 6002, 5878, 5757, 5640,
5527, 5417, 5310, 5207, 5106, 5008, 4913, 4820, 4731, 4643, 4558, 4475, 4395, 4317, 4240, 4166,
4093, 4023, 3954, 3887, 3821, 3758, 3696, 3635, 3576, 3518, 3462, 3407, 3352, 3300, 3250, 3200,
3151, 3103, 3056, 3010, 2966, 2922, 2879, 2837, 2796, 2756, 2717, 2679, 2641, 2604, 2568, 2533),
(163108, 162604, 161107, 158674, 155388, 151358, 146708, 141567, 136066, 130327, 124459, 118560, 112708, 106970, 101394, 96019,
90870, 85962, 81305, 76900, 72747, 68838, 65164, 61720, 58489, 55462, 52629, 49975, 47490, 45162, 42982, 40938,
39022, 37225, 35537, 33952, 32462, 31061, 29742, 28499, 27328, 26223, 25179, 24194, 23261, 22379, 21544, 20752,
20002, 19289, 18612, 17969, 17358, 16776, 16221, 15692, 15189, 14709, 14249, 13811, 13392, 12991, 12608, 12241,
11889, 11551, 11228, 10918, 10620, 10333, 10058, 9794, 9540, 9295, 9059, 8832, 8613, 8403, 8199, 8003,
7814, 7631, 7455, 7284, 7119, 6959, 6805, 6655, 6512, 6372, 6237, 6105, 5978, 5855, 5735, 5619,
5507, 5398, 5292, 5189, 5089, 4991, 4897, 4805, 4716, 4629, 4544, 4462, 4382, 4304, 4228, 4154,
4082, 4012, 3944, 3877, 3812, 3749, 3687, 3626, 3568, 3510, 3454, 3399, 3345, 3293, 3243, 3193,
3144, 3096, 3050, 3004, 2960, 2916, 2874, 2832, 2791, 2751, 2712, 2674, 2637, 2600, 2564, 2529),
(146391, 145984, 144777, 142809, 140142, 136855, 133042, 128801, 124231, 119429, 114484, 109473, 104465, 99517, 94674, 89971,
85434, 81082, 76926, 72972, 69221, 65673, 62322, 59163, 56188, 53390, 50759, 48285, 45962, 43778, 41726, 39798,
37984, 36279, 34675, 33164, 31741, 30400, 29135, 27942, 26815, 25750, 24743, 23791, 22889, 22034, 21224, 20455,
19725, 19032, 18373, 17746, 17149, 16581, 16039, 15522, 15029, 14559, 14109, 13679, 13268, 12874, 12498, 12137,
11791, 11459, 11140, 10835, 10541, 10259, 9988, 9727, 9476, 9235, 9002, 8778, 8562, 8353, 8151, 7958,
7771, 7591, 7416, 7247, 7084, 6926, 6773, 6625, 6482, 6344, 6209, 6079, 5953, 5831, 5712, 5597,
5486, 5377, 5272, 5170, 5071, 4974, 4880, 4789, 4700, 4614, 4530, 4448, 4369, 4291, 4216, 4142,
4071, 4000, 3932, 3867, 3802, 3739, 3676, 3617, 3558, 3502, 3445, 3391, 3338, 3286, 3234, 3186,
3137, 3090, 3043, 2998, 2954, 2910, 2868, 2826, 2786, 2746, 2707, 2669, 2632, 2595, 2559, 2524),
(132118, 131786, 130802, 129193, 127006, 124301, 121147, 117621, 113798, 109756, 105565, 101289, 96988, 92708, 88491, 84369,
80367, 76504, 72793, 69243, 65857, 62637, 59582, 56688, 53951, 51366, 48926, 46624, 44454, 42408, 40480, 38662,
36949, 35333, 33809, 32372, 31014, 29733, 28521, 27377, 26295, 25269, 24300, 23380, 22508, 21682, 20897, 20151,
19442, 18769, 18127, 17517, 16935, 16380, 15851, 15347, 14865, 14404, 13963, 13542, 13139, 12753, 12383, 12029,
11689, 11363, 11050, 10749, 10460, 10182, 9915, 9658, 9410, 9172, 8943, 8721, 8508, 8302, 8104, 7912,
7727, 7548, 7375, 7208, 7047, 6891, 6740, 6593, 6451, 6314, 6181, 6052, 5927, 5806, 5688, 5574,
5464, 5356, 5252, 5150, 5052, 4956, 4863, 4772, 4684, 4598, 4515, 4434, 4355, 4278, 4203, 4130,
4059, 3989, 3922, 3855, 3791, 3728, 3667, 3608, 3549, 3493, 3437, 3383, 3330, 3277, 3228, 3178,
3130, 3083, 3037, 2991, 2947, 2904, 2862, 2820, 2780, 2740, 2702, 2664, 2627, 2590, 2555, 2520),
(119835, 119561, 118751, 117424, 115614, 113369, 110739, 107785, 104567, 101143, 97574, 93910, 90201, 86488, 82806, 79186,
75650, 72218, 68902, 65713, 62656, 59734, 56949, 54300, 51784, 49397, 47137, 44996, 42972, 41057, 39247, 37536,
35919, 34390, 32945, 31579, 30286, 29062, 27904, 26808, 25768, 24784, 23850, 22964, 22122, 21323, 20563, 19841,
19154, 18499, 17876, 17282, 16715, 16175, 15659, 15165, 14695, 14245, 13814, 13402, 13007, 12628, 12266, 11918,
11584, 11263, 10956, 10660, 10376, 10102, 9839, 9586, 9342, 9107, 8881, 8663, 8452, 8249, 8053, 7864,
7681, 7504, 7334, 7167, 7009, 6854, 6704, 6560, 6419, 6283, 6152, 6024, 5900, 5780, 5663, 5550,
5441, 5334, 5230, 5130, 5032, 4937, 4844, 4755, 4667, 4582, 4499, 4419, 4340, 4264, 4189, 4117,
4046, 3977, 3910, 3844, 3780, 3718, 3657, 3598, 3540, 3483, 3428, 3374, 3321, 3270, 3220, 3170,
3122, 3075, 3029, 2984, 2941, 2898, 2855, 2814, 2774, 2735, 2696, 2658, 2621, 2585, 2549, 2515),
(109188, 108962, 108288, 107183, 105674, 103794, 101586, 99094, 96367, 93453, 90397, 87244, 84033, 80801, 77579, 74393,
71264, 68210, 65244, 62378, 59616, 56965, 54427, 52002, 49690, 47489, 45396, 43407, 41520, 39730, 38033, 36424,
34899, 33454, 32085, 30786, 29557, 28391, 27284, 26236, 25240, 24294, 23396, 22542, 21731, 20959, 20225, 19526,
18860, 18225, 17620, 17042, 16491, 15964, 15462, 14981, 14521, 14082, 13660, 13257, 12870, 12500, 12144, 11803,
11476, 11161, 10859, 10568, 10289, 10020, 9761, 9512, 9272, 9040, 8817, 8602, 8395, 8194, 8001, 7814,
7632, 7459, 7290, 7127, 6969, 6816, 6668, 6525, 6386, 6251, 6121, 5995, 5872, 5753, 5638, 5525,
5417, 5311, 5208, 5108, 5011, 4917, 4825, 4736, 4649, 4565, 4483, 4403, 4325, 4249, 4175, 4103,
4033, 3964, 3896, 3832, 3769, 3707, 3646, 3587, 3530, 3472, 3418, 3365, 3311, 3261, 3211, 3162,
3114, 3068, 3022, 2977, 2934, 2891, 2849, 2808, 2768, 2729, 2690, 2652, 2616, 2580, 2544, 2510),
(99900, 99710, 99146, 98219, 96950, 95366, 93498, 91384, 89059, 86564, 83936, 81211, 78422, 75600, 72772, 69961,
67187, 64466, 61810, 59231, 56736, 54330, 52015, 49797, 47673, 45643, 43706, 41860, 40102, 38430, 36840, 35328,
33892, 32528, 31232, 30001, 28832, 27721, 26665, 25662, 24709, 23802, 22939, 22118, 21336, 20592, 19882, 19206,
18562, 17946, 17359, 16798, 16263, 15751, 15261, 14793, 14344, 13915, 13503, 13109, 12731, 12368, 12020, 11686,
11365, 11056, 10759, 10474, 10199, 9935, 9681, 9435, 9199, 8971, 8752, 8540, 8335, 8137, 7947, 7761,
7584, 7412, 7245, 7084, 6927, 6777, 6630, 6489, 6351, 6218, 6089, 5964, 5843, 5725, 5611, 5500,
5392, 5287, 5185, 5086, 4990, 4897, 4806, 4717, 4631, 4547, 4466, 4386, 4309, 4234, 4160, 4089,
4018, 3951, 3884, 3820, 3757, 3694, 3635, 3576, 3519, 3463, 3409, 3355, 3302, 3252, 3202, 3154,
3106, 3060, 3014, 2970, 2926, 2884, 2842, 2801, 2761, 2722, 2684, 2647, 2610, 2574, 2539, 2504),
(91749, 91589, 91112, 90328, 89254, 87910, 86320, 84515, 82523, 80376, 78105, 75740, 73309, 70837, 68348, 65863,
63399, 60970, 58590, 56267, 54011, 51826, 49717, 47685, 45734, 43863, 42071, 40358, 38721, 37160, 35671, 34252,
32900, 31613, 30388, 29221, 28111, 27054, 26048, 25090, 24177, 23308, 22480, 21691, 20939, 20221, 19537, 18884,
18260, 17664, 17095, 16551, 16031, 15533, 15057, 14599, 14163, 13744, 13343, 12958, 12588, 12234, 11893, 11566,
11251, 10948, 10657, 10377, 10108, 9848, 9598, 9357, 9124, 8900, 8684, 8475, 8274, 8079, 7890, 7709,
7532, 7363, 7199, 7038, 6884, 6736, 6592, 6451, 6315, 6184, 6056, 5933, 5813, 5696, 5583, 5473,
5366, 5262, 5161, 5063, 4968, 4875, 4785, 4697, 4612, 4529, 4448, 4369, 4292, 4218, 4145, 4074,
4004, 3937, 3871, 3807, 3744, 3683, 3623, 3565, 3508, 3453, 3398, 3345, 3293, 3243, 3193, 3145,
3098, 3051, 3006, 2962, 2919, 2876, 2835, 2794, 2755, 2716, 2678, 2640, 2604, 2568, 2533, 2499),
(84555, 84420, 84014, 83348, 82432, 81284, 79924, 78373, 76658, 74802, 72831, 70770, 68643, 66471, 64275, 62072,
59879, 57708, 55571, 53477, 51435, 49450, 47526, 45666, 43874, 42148, 40491, 38902, 37379, 35922, 34529, 33198,
31926, 30713, 29554, 28449, 27397, 26392, 25433, 24519, 23647, 22815, 22021, 21264, 20540, 19849, 19189, 18559,
17956, 17380, 16828, 16300, 15795, 15312, 14849, 14405, 13980, 13572, 13180, 12803, 12443, 12096, 11763, 11443,
11135, 10838, 10553, 10278, 10014, 9759, 9513, 9276, 9048, 8827, 8615, 8409, 8211, 8019, 7833, 7654,
7481, 7313, 7151, 6994, 6841, 6694, 6551, 6413, 6279, 6149, 6023, 5900, 5781, 5666, 5554, 5445,
5339, 5237, 5137, 5040, 4945, 4853, 4764, 4677, 4592, 4510, 4430, 4352, 4275, 4201, 4129, 4058,
3990, 3923, 3857, 3793, 3731, 3670, 3611, 3553, 3497, 3442, 3388, 3334, 3283, 3232, 3184, 3136,
3089, 3043, 2998, 2954, 2911, 2869, 2827, 2787, 2748, 2709, 2671, 2634, 2598, 2562, 2527, 2493),
(78176, 78060, 77714, 77143, 76358, 75372, 74200, 72862, 71377, 69765, 68048, 66246, 64378, 62464, 60521, 58564,
56608, 54662, 52742, 50853, 49003, 47197, 45442, 43739, 42091, 40501, 38969, 37494, 36078, 34719, 33415, 32167,
30972, 29829, 28735, 27689, 26690, 25735, 24824, 23952, 23120, 22324, 21563, 20836, 20141, 19476, 18840, 18232,
17650, 17093, 16560, 16049, 15559, 15090, 14640, 14208, 13794, 13396, 13014, 12648, 12296, 11957, 11631, 11318,
11016, 10726, 10447, 10178, 9918, 9668, 9427, 9194, 8970, 8753, 8544, 8341, 8146, 7957, 7775, 7598,
7427, 7262, 7102, 6947, 6797, 6651, 6510, 6374, 6241, 6113, 5988, 5867, 5749, 5635, 5524, 5417,
5312, 5210, 5111, 5015, 4922, 4831, 4742, 4656, 4572, 4491, 4411, 4333, 4258, 4184, 4113, 4043,
3973, 3907, 3843, 3780, 3718, 3657, 3599, 3540, 3485, 3429, 3377, 3324, 3273, 3223, 3173, 3126,
3080, 3034, 2989, 2945, 2903, 2861, 2820, 2780, 2740, 2702, 2664, 2627, 2591, 2556, 2521, 2487),
(72493, 72393, 72095, 71603, 70926, 70075, 69061, 67901, 66609, 65203, 63701, 62119, 60474, 58782, 57058, 55315,
53567, 51822, 50093, 48385, 46707, 45064, 43461, 41901, 40387, 38920, 37503, 36135, 34818, 33550, 32332, 31162,
30039, 28962, 27931, 26942, 25995, 25089, 24221, 23391, 22596, 21835, 21107, 20409, 19742, 19103, 18491, 17905,
17343, 16805, 16289, 15794, 15320, 14865, 14428, 14008, 13605, 13219, 12847, 12489, 12146, 11815, 11497, 11191,
10896, 10612, 10338, 10075, 9820, 9575, 9338, 9110, 8890, 8677, 8471, 8272, 8080, 7894, 7715, 7541,
7371, 7209, 7052, 6899, 6751, 6607, 6468, 6333, 6202, 6075, 5952, 5833, 5716, 5604, 5494, 5387,
5284, 5183, 5085, 4990, 4898, 4808, 4720, 4634, 4551, 4470, 4392, 4315, 4240, 4167, 4096, 4025,
3959, 3893, 3828, 3765, 3703, 3644, 3586, 3529, 3472, 3418, 3365, 3313, 3262, 3213, 3164, 3117,
3070, 3025, 2980, 2937, 2894, 2853, 2812, 2772, 2733, 2694, 2657, 2620, 2584, 2549, 2515, 2481),
(67407, 67321, 67063, 66637, 66051, 65312, 64430, 63419, 62291, 61060, 59740, 58347, 56893, 55393, 53860, 52303,
50738, 49171, 47611, 46066, 44542, 43045, 41580, 40150, 38757, 37405, 36094, 34826, 33600, 32418, 31279, 30183,
29128, 28115, 27142, 26207, 25311, 24450, 23626, 22835, 22077, 21350, 20653, 19985, 19345, 18731, 18142, 17577,
17036, 16516, 16017, 15539, 15079, 14638, 14213, 13807, 13416, 13039, 12677, 12329, 11994, 11672, 11361, 11062,
10774, 10496, 10228, 9970, 9721, 9481, 9249, 9025, 8808, 8599, 8397, 8202, 8013, 7829, 7653, 7482,
7316, 7156, 7000, 6850, 6704, 6562, 6425, 6292, 6163, 6037, 5915, 5797, 5683, 5571, 5463, 5357,
5255, 5155, 5059, 4964, 4873, 4784, 4697, 4612, 4530, 4450, 4372, 4295, 4221, 4149, 4077, 4009,
3941, 3877, 3812, 3751, 3690, 3630, 3572, 3515, 3460, 3406, 3352, 3302, 3250, 3202, 3154, 3106,
3060, 3015, 2971, 2928, 2885, 2844, 2804, 2764, 2725, 2687, 2650, 2613, 2577, 2542, 2508, 2474),
(62838, 62763, 62539, 62169, 61658, 61014, 60244, 59358, 58369, 57287, 56123, 54891, 53603, 52270, 50903, 49511,
48105, 46694, 45285, 43885, 42500, 41136, 39795, 38483, 37202, 35954, 34742, 33565, 32425, 31323, 30259, 29231,
28241, 27287, 26370, 25487, 24638, 23822, 23039, 22286, 21563, 20869, 20203, 19563, 18949, 18360, 17794, 17250,
16728, 16227, 15745, 15283, 14838, 14410, 14000, 13604, 13224, 12858, 12506, 12167, 11841, 11527, 11224, 10932,
10650, 10379, 10117, 9864, 9620, 9385, 9157, 8938, 8725, 8520, 8322, 8130, 7944, 7764, 7589, 7421,
7259, 7101, 6948, 6798, 6655, 6516, 6381, 6249, 6122, 5998, 5878, 5761, 5648, 5538, 5431, 5327,
5225, 5127, 5031, 4938, 4847, 4759, 4673, 4589, 4508, 4428, 4351, 4276, 4202, 4130, 4059, 3991,
3926, 3861, 3796, 3735, 3675, 3615, 3558, 3502, 3447, 3394, 3341, 3290, 3240, 3191, 3143, 3096,
3050, 3005, 2962, 2919, 2877, 2835, 2795, 2756, 2717, 2679, 2642, 2606, 2570, 2535, 2501, 2468),
(58719, 58653, 58458, 58134, 57687, 57123, 56447, 55670, 54798, 53843, 52815, 51723, 50577, 49388, 48165, 46918,
45653, 44381, 43106, 41835, 40575, 39329, 38103, 36898, 35719, 34567, 33444, 32353, 31293, 30264, 29270, 28307,
27378, 26481, 25616, 24782, 23978, 23205, 22461, 21745, 21056, 20394, 19757, 19145, 18557, 17991, 17447, 16924,
16422, 15938, 15473, 15026, 14596, 14182, 13783, 13400, 13032, 12676, 12334, 12004, 11686, 11380, 11085, 10800,
10525, 10260, 10004, 9757, 9518, 9287, 9065, 8849, 8641, 8440, 8245, 8057, 7874, 7698, 7527, 7360,
7201, 7045, 6894, 6748, 6605, 6469, 6336, 6206, 6080, 5958, 5840, 5724, 5613, 5504, 5398, 5295,
5195, 5098, 5003, 4911, 4821, 4734, 4649, 4566, 4485, 4407, 4330, 4255, 4182, 4111, 4041, 3973,
3909, 3844, 3781, 3719, 3660, 3602, 3545, 3488, 3434, 3381, 3329, 3277, 3228, 3180, 3132, 3085,
3040, 2995, 2952, 2909, 2867, 2826, 2786, 2747, 2709, 2671, 2634, 2598, 2563, 2528, 2494, 2461),
(54992, 54934, 54762, 54478, 54086, 53589, 52994, 52308, 51537, 50693, 49780, 48809, 47787, 46725, 45629, 44507,
43368, 42218, 41063, 39908, 38760, 37622, 36497, 35391, 34304, 33241, 32201, 31188, 30202, 29243, 28313, 27411,
26539, 25695, 24880, 24092, 23333, 22600, 21893, 21212, 20557, 19925, 19317, 18731, 18168, 17625, 17103, 16600,
16116, 15650, 15201, 14770, 14354, 13954, 13568, 13197, 12839, 12494, 12161, 11840, 11531, 11233, 10945, 10667,
10399, 10140, 9890, 9648, 9415, 9189, 8971, 8760, 8556, 8358, 8167, 7982, 7803, 7630, 7462, 7299,
7141, 6988, 6840, 6696, 6555, 6421, 6290, 6162, 6038, 5918, 5801, 5687, 5576, 5469, 5365, 5263,
5164, 5068, 4974, 4883, 4795, 4708, 4624, 4542, 4462, 4384, 4308, 4234, 4162, 4092, 4023, 3956,
3891, 3827, 3765, 3703, 3645, 3587, 3530, 3475, 3420, 3368, 3316, 3266, 3216, 3168, 3121, 3074,
3029, 2985, 2942, 2899, 2858, 2817, 2777, 2739, 2700, 2663, 2626, 2590, 2555, 2521, 2487, 2454),
(51609, 51558, 51405, 51156, 50810, 50371, 49845, 49238, 48555, 47804, 46991, 46125, 45212, 44259, 43275, 42265,
41236, 40195, 39146, 38096, 37048, 36007, 34976, 33958, 32957, 31974, 31011, 30070, 29152, 28258, 27389, 26544,
25724, 24932, 24163, 23420, 22701, 22007, 21336, 20689, 20065, 19463, 18882, 18322, 17782, 17262, 16761, 16278,
15812, 15364, 14931, 14515, 14113, 13726, 13352, 12992, 12645, 12310, 11987, 11675, 11375, 11084, 10804, 10533,
10271, 10019, 9774, 9538, 9310, 9089, 8876, 8669, 8469, 8276, 8089, 7907, 7731, 7561, 7396, 7235,
7081, 6931, 6784, 6643, 6506, 6372, 6243, 6117, 5995, 5876, 5761, 5649, 5540, 5434, 5330, 5230,
5133, 5038, 4945, 4855, 4767, 4682, 4599, 4518, 4439, 4362, 4286, 4213, 4142, 4072, 4004, 3938,
3873, 3810, 3748, 3688, 3629, 3571, 3515, 3460, 3407, 3354, 3302, 3253, 3204, 3156, 3109, 3063,
3018, 2974, 2931, 2889, 2848, 2808, 2768, 2730, 2692, 2655, 2618, 2583, 2548, 2513, 2480, 2447),
(48528, 48483, 48349, 48128, 47821, 47433, 46966, 46426, 45819, 45149, 44424, 43649, 42830, 41974, 41088, 40176,
39246, 38301, 37348, 36391, 35433, 34480, 33533, 32597, 31673, 30764, 29872, 28997, 28143, 27309, 26495, 25705,
24936, 24190, 23466, 22764, 22085, 21427, 20791, 20176, 19582, 19008, 18453, 17918, 17402, 16903, 16422, 15958,
15511, 15079, 14662, 14260, 13872, 13497, 13136, 12788, 12451, 12127, 11813, 11510, 11218, 10935, 10662, 10398,
10143, 9897, 9658, 9428, 9205, 8989, 8780, 8578, 8382, 8192, 8008, 7831, 7659, 7491, 7328, 7172,
7020, 6872, 6728, 6589, 6454, 6322, 6195, 6071, 5951, 5834, 5720, 5610, 5502, 5397, 5296, 5197,
5100, 5006, 4915, 4826, 4740, 4655, 4573, 4493, 4414, 4338, 4264, 4191, 4121, 4052, 3984, 3919,
3855, 3792, 3731, 3671, 3613, 3556, 3500, 3445, 3393, 3341, 3290, 3240, 3191, 3144, 3097, 3052,
3007, 2964, 2921, 2879, 2838, 2798, 2759, 2720, 2683, 2646, 2610, 2574, 2540, 2506, 2472, 2439),
(45716, 45676, 45557, 45360, 45088, 44742, 44327, 43846, 43303, 42705, 42055, 41360, 40624, 39853, 39053, 38229,
37386, 36528, 35660, 34786, 33910, 33036, 32166, 31302, 30450, 29609, 28782, 27969, 27173, 26395, 25635, 24894,
24172, 23470, 22788, 22126, 21483, 20860, 20257, 19673, 19107, 18560, 18032, 17520, 17026, 16549, 16087, 15642,
15212, 14796, 14395, 14007, 13632, 13271, 12921, 12584, 12258, 11943, 11639, 11345, 11060, 10786, 10520, 10263,
10014, 9774, 9541, 9316, 9098, 8888, 8683, 8486, 8294, 8108, 7928, 7754, 7585, 7421, 7262, 7108,
6958, 6813, 6672, 6535, 6401, 6272, 6147, 6025, 5906, 5791, 5679, 5570, 5464, 5361, 5260, 5163,
5068, 4975, 4885, 4797, 4711, 4628, 4546, 4467, 4390, 4315, 4241, 4169, 4099, 4031, 3964, 3898,
3836, 3774, 3713, 3654, 3596, 3540, 3485, 3431, 3377, 3326, 3275, 3227, 3179, 3130, 3085, 3040,
2996, 2953, 2910, 2869, 2828, 2788, 2749, 2711, 2674, 2637, 2601, 2566, 2531, 2498, 2464, 2432),
(43141, 43105, 42999, 42824, 42581, 42273, 41902, 41471, 40986, 40449, 39866, 39241, 38578, 37882, 37159, 36412,
35646, 34865, 34073, 33275, 32472, 31669, 30869, 30074, 29286, 28507, 27739, 26984, 26242, 25516, 24805, 24110,
23433, 22772, 22129, 21504, 20897, 20307, 19735, 19180, 18642, 18121, 17617, 17128, 16656, 16199, 15756, 15329,
14915, 14516, 14129, 13755, 13394, 13045, 12706, 12381, 12065, 11760, 11464, 11179, 10903, 10636, 10377, 10127,
9885, 9651, 9424, 9204, 8992, 8786, 8586, 8393, 8205, 8023, 7847, 7675, 7510, 7350, 7194, 7042,
6895, 6753, 6614, 6479, 6349, 6221, 6098, 5978, 5861, 5748, 5637, 5530, 5425, 5324, 5225, 5128,
5034, 4943, 4854, 4767, 4682, 4600, 4520, 4441, 4365, 4290, 4218, 4147, 4077, 4009, 3944, 3880,
3817, 3755, 3694, 3637, 3580, 3524, 3469, 3415, 3363, 3311, 3262, 3213, 3164, 3119, 3073, 3028,
2984, 2941, 2899, 2858, 2818, 2778, 2739, 2702, 2664, 2628, 2592, 2557, 2523, 2490, 2457, 2424),
(40777, 40745, 40651, 40494, 40277, 40001, 39668, 39283, 38847, 38365, 37839, 37276, 36677, 36048, 35392, 34713,
34017, 33305, 32582, 31851, 31115, 30377, 29640, 28906, 28177, 27455, 26743, 26040, 25349, 24670, 24005, 23354,
22717, 22096, 21491, 20900, 20326, 19768, 19225, 18698, 18187, 17691, 17209, 16743, 16291, 15853, 15430, 15020,
14621, 14238, 13866, 13506, 13157, 12820, 12494, 12178, 11872, 11577, 11291, 11014, 10745, 10486, 10235, 9991,
9756, 9527, 9306, 9092, 8884, 8683, 8488, 8299, 8116, 7938, 7765, 7598, 7435, 7278, 7124, 6976,
6832, 6691, 6555, 6422, 6295, 6170, 6048, 5930, 5815, 5704, 5595, 5489, 5386, 5286, 5188, 5093,
5000, 4910, 4822, 4737, 4653, 4572, 4492, 4415, 4339, 4266, 4194, 4124, 4055, 3988, 3923, 3860,
3796, 3737, 3676, 3619, 3562, 3506, 3453, 3400, 3348, 3297, 3248, 3198, 3152, 3106, 3060, 3016,
2972, 2930, 2888, 2847, 2807, 2768, 2729, 2692, 2655, 2619, 2583, 2549, 2515, 2481, 2448, 2416),
(38603, 38574, 38490, 38349, 38154, 37906, 37608, 37261, 36869, 36434, 35960, 35450, 34908, 34338, 33742, 33125,
32490, 31840, 31178, 30508, 29833, 29154, 28474, 27796, 27121, 26451, 25790, 25135, 24491, 23857, 23234, 22624,
22026, 21442, 20871, 20314, 19771, 19242, 18728, 18227, 17741, 17269, 16810, 16364, 15933, 15514, 15108, 14714,
14333, 13963, 13605, 13258, 12922, 12597, 12282, 11977, 11681, 11395, 11117, 10849, 10588, 10336, 10092, 9855,
9626, 9404, 9188, 8979, 8777, 8580, 8390, 8205, 8026, 7852, 7683, 7519, 7360, 7205, 7055, 6909,
6768, 6630, 6497, 6367, 6241, 6118, 5998, 5882, 5769, 5659, 5552, 5448, 5346, 5247, 5151, 5057,
4966, 4877, 4790, 4706, 4623, 4543, 4465, 4388, 4314, 4241, 4170, 4100, 4033, 3966, 3902, 3839,
3778, 3717, 3658, 3601, 3545, 3490, 3436, 3384, 3333, 3282, 3232, 3185, 3138, 3092, 3047, 3003,
2960, 2918, 2876, 2836, 2796, 2757, 2719, 2682, 2645, 2609, 2574, 2540, 2506, 2473, 2440, 2408),
(36598, 36572, 36496, 36370, 36194, 35971, 35702, 35389, 35035, 34643, 34214, 33752, 33261, 32742, 32200, 31638,
31058, 30463, 29857, 29242, 28621, 27994, 27367, 26740, 26116, 25495, 24879, 24270, 23668, 23076, 22493, 21920,
21359, 20809, 20271, 19745, 19231, 18731, 18243, 17768, 17305, 16855, 16418, 15992, 15580, 15179, 14791, 14413,
14047, 13691, 13347, 13013, 12690, 12376, 12071, 11776, 11490, 11213, 10945, 10684, 10432, 10187, 9949, 9719,
9496, 9280, 9070, 8866, 8669, 8477, 8291, 8110, 7935, 7765, 7600, 7439, 7284, 7131, 6984, 6843,
6704, 6569, 6438, 6310, 6186, 6065, 5948, 5833, 5722, 5614, 5509, 5406, 5306, 5209, 5114, 5021,
4931, 4844, 4758, 4675, 4593, 4514, 4437, 4361, 4287, 4215, 4145, 4077, 4009, 3944, 3880, 3818,
3757, 3698, 3640, 3583, 3527, 3472, 3420, 3368, 3317, 3266, 3219, 3171, 3124, 3079, 3034, 2990,
2948, 2906, 2865, 2824, 2785, 2747, 2709, 2672, 2635, 2600, 2565, 2531, 2497, 2464, 2432, 2400),
(34745, 34722, 34653, 34539, 34381, 34180, 33937, 33654, 33334, 32978, 32589, 32170, 31723, 31251, 30757, 30244,
29713, 29169, 28613, 28047, 27475, 26898, 26318, 25738, 25158, 24582, 24009, 23441, 22879, 22325, 21779, 21242,
20714, 20196, 19689, 19193, 18707, 18233, 17771, 17319, 16880, 16451, 16035, 15629, 15235, 14851, 14479, 14116,
13765, 13424, 13092, 12770, 12459, 12157, 11863, 11578, 11301, 11033, 10773, 10520, 10275, 10038, 9807, 9584,
9367, 9156, 8951, 8753, 8561, 8374, 8192, 8015, 7845, 7678, 7517, 7360, 7206, 7059, 6915, 6775,
6639, 6506, 6378, 6252, 6131, 6012, 5897, 5784, 5675, 5568, 5465, 5364, 5265, 5169, 5076, 4985,
4896, 4810, 4725, 4643, 4563, 4484, 4408, 4333, 4261, 4190, 4120, 4052, 3986, 3922, 3859, 3796,
3737, 3678, 3620, 3564, 3509, 3454, 3403, 3351, 3300, 3252, 3204, 3156, 3110, 3065, 3021, 2977,
2935, 2893, 2853, 2813, 2774, 2736, 2698, 2661, 2625, 2590, 2555, 2521, 2488, 2455, 2423, 2392),
(33029, 33009, 32947, 32844, 32700, 32518, 32298, 32042, 31752, 31429, 31075, 30694, 30286, 29857, 29404, 28935,
28449, 27950, 27439, 26919, 26390, 25857, 25322, 24785, 24247, 23711, 23177, 22647, 22123, 21604, 21092, 20588,
20092, 19604, 19126, 18657, 18198, 17749, 17311, 16882, 16464, 16056, 15659, 15272, 14895, 14529, 14172, 13825,
13488, 13160, 12842, 12531, 12231, 11940, 11656, 11381, 11113, 10854, 10602, 10357, 10120, 9889, 9666, 9448,
9237, 9032, 8833, 8640, 8452, 8270, 8093, 7921, 7754, 7591, 7432, 7280, 7130, 6984, 6844, 6707,
6574, 6444, 6317, 6195, 6075, 5958, 5845, 5735, 5627, 5522, 5420, 5321, 5224, 5130, 5038, 4948,
4861, 4775, 4692, 4611, 4532, 4455, 4379, 4306, 4234, 4164, 4095, 4028, 3963, 3898, 3837, 3776,
3716, 3658, 3601, 3545, 3490, 3438, 3386, 3334, 3284, 3236, 3188, 3141, 3096, 3051, 3007, 2964,
2922, 2881, 2841, 2801, 2762, 2724, 2687, 2651, 2615, 2580, 2546, 2512, 2479, 2446, 2414, 2383),
(31438, 31419, 31363, 31269, 31140, 30974, 30775, 30542, 30278, 29984, 29663, 29315, 28943, 28549, 28137, 27707,
27261, 26801, 26332, 25852, 25365, 24873, 24376, 23878, 23378, 22879, 22382, 21888, 21397, 20912, 20432, 19958,
19492, 19032, 18581, 18139, 17705, 17279, 16863, 16456, 16059, 15670, 15292, 14923, 14563, 14212, 13871, 13538,
13214, 12900, 12594, 12296, 12006, 11725, 11451, 11186, 10927, 10676, 10432, 10196, 9965, 9742, 9524, 9313,
9108, 8909, 8715, 8527, 8344, 8167, 7994, 7826, 7663, 7504, 7349, 7199, 7053, 6911, 6773, 6639,
6508, 6381, 6257, 6136, 6019, 5904, 5793, 5685, 5579, 5476, 5376, 5278, 5183, 5090, 4999, 4911,
4825, 4741, 4659, 4579, 4501, 4424, 4350, 4277, 4206, 4137, 4070, 4003, 3939, 3876, 3814, 3753,
3694, 3638, 3581, 3526, 3472, 3420, 3368, 3318, 3268, 3220, 3173, 3127, 3081, 3037, 2993, 2951,
2909, 2868, 2828, 2789, 2751, 2713, 2676, 2640, 2605, 2570, 2536, 2502, 2469, 2437, 2406, 2375),
(29959, 29942, 29891, 29806, 29687, 29537, 29356, 29143, 28904, 28636, 28342, 28025, 27685, 27325, 26945, 26551,
26142, 25718, 25285, 24843, 24393, 23938, 23478, 23015, 22550, 22086, 21622, 21160, 20702, 20247, 19796, 19352,
18913, 18480, 18054, 17636, 17226, 16823, 16428, 16042, 15664, 15294, 14934, 14581, 14237, 13902, 13575, 13256,
12946, 12644, 12349, 12063, 11784, 11513, 11249, 10993, 10743, 10500, 10264, 10035, 9812, 9595, 9384, 9179,
8980, 8786, 8598, 8414, 8236, 8062, 7895, 7731, 7571, 7416, 7266, 7119, 6976, 6837, 6702, 6569,
6442, 6317, 6196, 6078, 5962, 5850, 5741, 5634, 5531, 5429, 5331, 5235, 5141, 5049, 4960, 4873,
4788, 4706, 4625, 4546, 4469, 4394, 4320, 4249, 4179, 4110, 4043, 3978, 3914, 3852, 3792, 3732,
3674, 3617, 3561, 3506, 3453, 3401, 3350, 3300, 3252, 3204, 3157, 3111, 3066, 3022, 2979, 2937,
2896, 2856, 2816, 2777, 2739, 2702, 2665, 2629, 2594, 2559, 2526, 2492, 2460, 2428, 2397, 2366),
(28581, 28566, 28519, 28442, 28335, 28198, 28032, 27839, 27620, 27375, 27106, 26816, 26505, 26173, 25827, 25463,
25087, 24698, 24298, 23889, 23472, 23050, 22623, 22193, 21761, 21328, 20895, 20464, 20034, 19608, 19186, 18767,
18354, 17947, 17545, 17150, 16761, 16380, 16005, 15638, 15279, 14927, 14582, 14247, 13919, 13597, 13285, 12980,
12681, 12392, 12109, 11833, 11565, 11304, 11049, 10802, 10560, 10326, 10098, 9875, 9659, 9449, 9245, 9046,
8852, 8664, 8480, 8302, 8129, 7960, 7796, 7636, 7480, 7328, 7181, 7038, 6899, 6763, 6630, 6501,
6376, 6254, 6135, 6019, 5906, 5796, 5688, 5584, 5482, 5382, 5285, 5191, 5099, 5009, 4921, 4835,
4752, 4670, 4591, 4513, 4437, 4363, 4291, 4220, 4151, 4083, 4018, 3953, 3889, 3828, 3769, 3710,
3651, 3596, 3540, 3487, 3434, 3383, 3332, 3283, 3234, 3187, 3141, 3096, 3051, 3008, 2965, 2923,
2883, 2842, 2803, 2765, 2727, 2690, 2654, 2618, 2583, 2549, 2515, 2482, 2450, 2418, 2387, 2357),
(27297, 27283, 27239, 27170, 27072, 26947, 26795, 26619, 26418, 26194, 25949, 25682, 25396, 25093, 24774, 24439,
24092, 23733, 23363, 22985, 22599, 22207, 21811, 21411, 21008, 20605, 20200, 19797, 19395, 18995, 18598, 18205,
17816, 17432, 17052, 16679, 16311, 15950, 15594, 15246, 14904, 14568, 14241, 13921, 13607, 13300, 13000, 12708,
12423, 12144, 11872, 11607, 11349, 11097, 10852, 10613, 10380, 10153, 9932, 9717, 9508, 9304, 9106, 8913,
8725, 8542, 8364, 8190, 8021, 7857, 7697, 7541, 7389, 7242, 7098, 6958, 6821, 6687, 6559, 6433,
6310, 6190, 6074, 5960, 5849, 5741, 5636, 5533, 5433, 5335, 5240, 5147, 5056, 4968, 4881, 4797,
4715, 4635, 4556, 4480, 4405, 4332, 4261, 4191, 4123, 4056, 3991, 3928, 3864, 3805, 3744, 3687,
3630, 3574, 3520, 3467, 3415, 3364, 3314, 3265, 3218, 3171, 3125, 3080, 3036, 2993, 2951, 2909,
2869, 2829, 2790, 2752, 2715, 2678, 2642, 2607, 2572, 2538, 2505, 2472, 2440, 2409, 2378, 2348),
(26096, 26084, 26046, 25981, 25892, 25777, 25639, 25477, 25293, 25088, 24862, 24617, 24355, 24076, 23781, 23473,
23152, 22821, 22479, 22128, 21771, 21407, 21038, 20666, 20290, 19914, 19536, 19158, 18781, 18406, 18033, 17663,
17297, 16934, 16576, 16223, 15875, 15532, 15195, 14864, 14539, 14220, 13908, 13602, 13302, 13009, 12722, 12442,
12168, 11901, 11639, 11385, 11136, 10894, 10657, 10426, 10202, 9983, 9769, 9561, 9358, 9161, 8968, 8781,
8598, 8421, 8247, 8079, 7914, 7754, 7598, 7446, 7299, 7154, 7013, 6877, 6744, 6614, 6487, 6364,
6244, 6126, 6012, 5901, 5792, 5686, 5583, 5482, 5383, 5288, 5194, 5103, 5014, 4927, 4842, 4759,
4678, 4599, 4522, 4446, 4372, 4301, 4230, 4161, 4093, 4029, 3965, 3902, 3839, 3780, 3722, 3664,
3608, 3553, 3500, 3447, 3395, 3345, 3296, 3248, 3200, 3154, 3109, 3064, 3021, 2978, 2936, 2895,
2855, 2816, 2777, 2739, 2702, 2666, 2630, 2595, 2561, 2527, 2494, 2462, 2430, 2399, 2368, 2338),
(24975, 24963, 24928, 24869, 24786, 24682, 24555, 24406, 24237, 24049, 23841, 23616, 23375, 23117, 22846, 22561,
22265, 21958, 21641, 21316, 20984, 20646, 20303, 19956, 19605, 19253, 18900, 18546, 18193, 17841, 17490, 17142,
16797, 16455, 16116, 15781, 15453, 15128, 14807, 14493, 14184, 13880, 13583, 13289, 13003, 12724, 12449, 12181,
11918, 11662, 11411, 11166, 10927, 10693, 10465, 10243, 10026, 9814, 9607, 9406, 9210, 9019, 8832, 8650,
8473, 8300, 8132, 7968, 7808, 7652, 7500, 7352, 7208, 7067, 6930, 6797, 6666, 6539, 6415, 6295,
6177, 6062, 5950, 5841, 5735, 5631, 5529, 5431, 5334, 5240, 5148, 5058, 4971, 4885, 4802, 4720,
4640, 4563, 4487, 4412, 4340, 4269, 4200, 4132, 4066, 4000, 3938, 3876, 3815, 3756, 3698, 3641,
3586, 3531, 3479, 3427, 3376, 3326, 3277, 3229, 3182, 3137, 3092, 3048, 3005, 2963, 2921, 2881,
2841, 2802, 2764, 2727, 2690, 2654, 2619, 2584, 2550, 2517, 2484, 2452, 2420, 2389, 2359, 2329),
(23924, 23913, 23880, 23826, 23750, 23654, 23538, 23401, 23246, 23072, 22881, 22674, 22451, 22214, 21963, 21700,
21425, 21141, 20847, 20545, 20237, 19922, 19602, 19279, 18952, 18622, 18292, 17960, 17629, 17298, 16968, 16640,
16314, 15992, 15672, 15356, 15043, 14735, 14432, 14133, 13839, 13549, 13264, 12987, 12713, 12445, 12182, 11925,
11673, 11427, 11186, 10951, 10720, 10495, 10276, 10061, 9852, 9647, 9448, 9253, 9063, 8878, 8697, 8521,
8349, 8180, 8017, 7858, 7702, 7550, 7403, 7258, 7117, 6980, 6847, 6716, 6589, 6465, 6344, 6226,
6111, 5998, 5889, 5782, 5677, 5576, 5476, 5379, 5284, 5192, 5102, 5014, 4928, 4843, 4761, 4681,
4603, 4526, 4451, 4378, 4307, 4237, 4169, 4102, 4037, 3973, 3911, 3850, 3790, 3731, 3674, 3617,
3564, 3510, 3458, 3406, 3356, 3307, 3258, 3211, 3164, 3120, 3075, 3032, 2989, 2947, 2906, 2866,
2827, 2788, 2751, 2714, 2677, 2641, 2606, 2572, 2538, 2505, 2473, 2441, 2410, 2379, 2349, 2320),
(22937, 22927, 22897, 22847, 22778, 22689, 22582, 22457, 22314, 22154, 21977, 21786, 21580, 21361, 21129, 20885,
20631, 20367, 20094, 19814, 19526, 19233, 18935, 18633, 18327, 18019, 17709, 17398, 17087, 16776, 16466, 16157,
15850, 15545, 15242, 14943, 14646, 14355, 14066, 13783, 13503, 13227, 12956, 12690, 12429, 12173, 11921, 11675,
11433, 11197, 10966, 10739, 10518, 10301, 10089, 9882, 9680, 9483, 9290, 9102, 8918, 8738, 8563, 8392,
8225, 8062, 7903, 7747, 7597, 7449, 7305, 7165, 7027, 6894, 6763, 6636, 6512, 6390, 6272, 6157,
6044, 5934, 5827, 5722, 5620, 5520, 5423, 5328, 5235, 5144, 5055, 4969, 4884, 4802, 4721, 4642,
4565, 4490, 4416, 4344, 4274, 4205, 4138, 4072, 4007, 3945, 3883, 3823, 3764, 3707, 3649, 3595,
3540, 3488, 3436, 3385, 3336, 3287, 3239, 3193, 3147, 3102, 3058, 3015, 2973, 2932, 2891, 2852,
2813, 2775, 2737, 2700, 2664, 2629, 2594, 2560, 2527, 2494, 2462, 2430, 2399, 2369, 2339, 2310),
(22010, 22001, 21974, 21928, 21864, 21782, 21683, 21568, 21436, 21288, 21125, 20948, 20758, 20555, 20340, 20114,
19878, 19633, 19379, 19118, 18851, 18577, 18299, 18017, 17731, 17442, 17152, 16860, 16567, 16275, 15983, 15691,
15401, 15114, 14828, 14544, 14263, 13987, 13713, 13443, 13175, 12914, 12656, 12402, 12152, 11907, 11666, 11430,
11198, 10972, 10749, 10532, 10319, 10110, 9906, 9706, 9511, 9321, 9134, 8952, 8774, 8600, 8430, 8265,
8103, 7945, 7790, 7640, 7492, 7349, 7209, 7072, 6938, 6808, 6680, 6555, 6435, 6317, 6201, 6088,
5978, 5870, 5765, 5663, 5563, 5465, 5369, 5276, 5185, 5096, 5009, 4924, 4841, 4760, 4680, 4603,
4527, 4453, 4381, 4310, 4241, 4173, 4107, 4041, 3978, 3916, 3855, 3796, 3737, 3681, 3626, 3571,
3518, 3466, 3415, 3365, 3315, 3266, 3220, 3173, 3129, 3085, 3041, 2999, 2957, 2916, 2876, 2837,
2798, 2760, 2723, 2687, 2651, 2616, 2582, 2548, 2515, 2483, 2451, 2420, 2389, 2359, 2329, 2300),
(21139, 21130, 21105, 21063, 21004, 20928, 20837, 20730, 20608, 20472, 20321, 20157, 19981, 19793, 19593, 19384,
19164, 18936, 18700, 18457, 18208, 17953, 17693, 17428, 17161, 16890, 16618, 16344, 16069, 15792, 15518, 15243,
14970, 14696, 14427, 14159, 13893, 13630, 13369, 13111, 12859, 12609, 12362, 12120, 11881, 11647, 11417, 11190,
10968, 10751, 10537, 10328, 10123, 9922, 9725, 9533, 9345, 9161, 8981, 8804, 8632, 8464, 8299, 8139,
7982, 7828, 7678, 7532, 7389, 7249, 7113, 6979, 6848, 6722, 6598, 6476, 6358, 6243, 6130, 6020,
5912, 5807, 5704, 5603, 5505, 5409, 5316, 5224, 5135, 5048, 4962, 4879, 4797, 4718, 4640, 4564,
4489, 4416, 4345, 4275, 4207, 4140, 4075, 4011, 3948, 3888, 3828, 3769, 3712, 3656, 3601, 3547,
3495, 3443, 3393, 3343, 3295, 3248, 3200, 3155, 3111, 3067, 3024, 2982, 2941, 2900, 2861, 2822,
2784, 2746, 2710, 2674, 2638, 2604, 2570, 2536, 2503, 2471, 2440, 2409, 2378, 2348, 2319, 2290),
(20318, 20310, 20287, 20248, 20193, 20123, 20039, 19940, 19827, 19701, 19561, 19410, 19246, 19071, 18886, 18691,
18487, 18275, 18055, 17828, 17595, 17357, 17114, 16867, 16616, 16361, 16106, 15849, 15590, 15331, 15071, 14812,
14553, 14296, 14040, 13786, 13533, 13284, 13036, 12792, 12550, 12312, 12077, 11846, 11618, 11393, 11173, 10956,
10743, 10534, 10329, 10128, 9931, 9737, 9548, 9362, 9181, 9003, 8829, 8659, 8492, 8329, 8169, 8014,
7861, 7713, 7567, 7425, 7285, 7149, 7017, 6887, 6761, 6637, 6516, 6397, 6282, 6169, 6059, 5951,
5846, 5743, 5642, 5544, 5448, 5354, 5262, 5173, 5085, 4999, 4916, 4834, 4754, 4675, 4599, 4524,
4451, 4379, 4309, 4241, 4174, 4108, 4043, 3981, 3919, 3859, 3800, 3743, 3685, 3631, 3577, 3524,
3472, 3420, 3370, 3322, 3274, 3228, 3182, 3137, 3092, 3049, 3007, 2965, 2924, 2884, 2845, 2807,
2769, 2732, 2696, 2660, 2625, 2591, 2557, 2524, 2492, 2460, 2428, 2398, 2368, 2338, 2309, 2280),
(19544, 19537, 19515, 19479, 19428, 19364, 19286, 19194, 19089, 18972, 18843, 18702, 18550, 18388, 18216, 18034,
17844, 17646, 17441, 17230, 17012, 16789, 16561, 16330, 16095, 15856, 15616, 15373, 15129, 14886, 14641, 14396,
14152, 13908, 13666, 13425, 13186, 12948, 12713, 12481, 12251, 12024, 11799, 11578, 11360, 11146, 10935, 10727,
10523, 10322, 10125, 9932, 9742, 9556, 9374, 9195, 9019, 8848, 8680, 8515, 8354, 8196, 8042, 7890,
7743, 7599, 7457, 7319, 7184, 7052, 6923, 6796, 6673, 6551, 6433, 6319, 6206, 6096, 5988, 5883,
5780, 5679, 5581, 5485, 5391, 5299, 5209, 5121, 5035, 4951, 4869, 4789, 4710, 4633, 4558, 4485,
4413, 4342, 4273, 4206, 4140, 4075, 4012, 3950, 3889, 3830, 3771, 3716, 3660, 3605, 3552, 3500,
3447, 3398, 3349, 3300, 3254, 3207, 3162, 3117, 3074, 3031, 2989, 2948, 2908, 2868, 2829, 2791,
2754, 2717, 2682, 2646, 2612, 2578, 2544, 2512, 2480, 2448, 2417, 2387, 2357, 2327, 2299, 2270),
(18814, 18807, 18787, 18753, 18706, 18647, 18574, 18489, 18392, 18283, 18163, 18032, 17891, 17740, 17579, 17410,
17233, 17049, 16857, 16659, 16456, 16247, 16034, 15817, 15595, 15372, 15146, 14918, 14689, 14457, 14227, 13996,
13765, 13533, 13305, 13075, 12849, 12624, 12400, 12179, 11960, 11743, 11529, 11318, 11110, 10904, 10702, 10503,
10307, 10115, 9926, 9740, 9557, 9378, 9202, 9030, 8861, 8695, 8532, 8373, 8217, 8065, 7915, 7768,
7625, 7486, 7348, 7214, 7083, 6954, 6829, 6705, 6585, 6468, 6353, 6240, 6130, 6023, 5918, 5815,
5714, 5616, 5520, 5426, 5334, 5244, 5156, 5070, 4985, 4903, 4822, 4744, 4666, 4591, 4517, 4445,
4374, 4305, 4237, 4171, 4106, 4043, 3980, 3920, 3860, 3802, 3744, 3688, 3633, 3580, 3527, 3476,
3425, 3375, 3327, 3279, 3232, 3187, 3141, 3098, 3055, 3013, 2972, 2931, 2891, 2852, 2814, 2776,
2739, 2703, 2667, 2632, 2598, 2565, 2532, 2499, 2467, 2436, 2405, 2375, 2346, 2317, 2288, 2260),
(18123, 18117, 18098, 18067, 18024, 17968, 17901, 17822, 17732, 17630, 17519, 17397, 17265, 17125, 16975, 16818,
16652, 16480, 16300, 16116, 15925, 15730, 15530, 15326, 15118, 14907, 14695, 14481, 14263, 14047, 13829, 13610,
13392, 13173, 12956, 12739, 12523, 12309, 12096, 11886, 11677, 11470, 11266, 11064, 10865, 10669, 10475, 10284,
10097, 9912, 9730, 9551, 9376, 9203, 9034, 8868, 8705, 8544, 8388, 8234, 8083, 7935, 7790, 7649,
7510, 7374, 7241, 7110, 6983, 6858, 6734, 6616, 6499, 6383, 6272, 6163, 6055, 5950, 5848, 5747,
5649, 5553, 5459, 5367, 5277, 5189, 5102, 5018, 4936, 4855, 4776, 4698, 4623, 4549, 4476, 4405,
4336, 4268, 4201, 4136, 4072, 4009, 3948, 3889, 3830, 3771, 3716, 3660, 3607, 3554, 3502, 3451,
3401, 3352, 3305, 3258, 3212, 3166, 3122, 3079, 3036, 2995, 2954, 2914, 2874, 2836, 2798, 2761,
2724, 2688, 2653, 2618, 2585, 2551, 2519, 2487, 2455, 2424, 2394, 2364, 2335, 2306, 2278, 2250),
(17470, 17464, 17447, 17418, 17378, 17326, 17263, 17190, 17106, 17012, 16908, 16794, 16672, 16540, 16401, 16253,
16099, 15938, 15770, 15597, 15419, 15235, 15048, 14856, 14660, 14463, 14263, 14061, 13857, 13652, 13444, 13239,
13032, 12825, 12617, 12413, 12208, 12004, 11802, 11601, 11402, 11205, 11010, 10817, 10627, 10439, 10254, 10071,
9891, 9713, 9539, 9367, 9198, 9032, 8869, 8708, 8551, 8397, 8245, 8096, 7950, 7807, 7667, 7530,
7395, 7263, 7134, 7006, 6883, 6762, 6643, 6526, 6413, 6301, 6192, 6085, 5981, 5878, 5778, 5680,
5584, 5490, 5398, 5308, 5220, 5134, 5049, 4967, 4886, 4807, 4729, 4653, 4579, 4506, 4435, 4366,
4297, 4231, 4165, 4101, 4038, 3977, 3917, 3858, 3800, 3743, 3688, 3633, 3580, 3528, 3477, 3427,
3377, 3330, 3282, 3236, 3191, 3146, 3102, 3060, 3018, 2976, 2936, 2896, 2857, 2819, 2782, 2745,
2709, 2673, 2639, 2604, 2571, 2538, 2506, 2474, 2443, 2412, 2382, 2352, 2323, 2295, 2267, 2239),
(16852, 16846, 16830, 16803, 16766, 16718, 16659, 16591, 16513, 16425, 16328, 16222, 16108, 15985, 15855, 15717,
15573, 15422, 15265, 15103, 14935, 14763, 14587, 14407, 14223, 14037, 13848, 13657, 13465, 13271, 13075, 12880,
12684, 12488, 12293, 12097, 11903, 11709, 11516, 11325, 11136, 10948, 10761, 10577, 10395, 10215, 10037, 9862,
9689, 9519, 9351, 9186, 9024, 8864, 8706, 8552, 8400, 8251, 8105, 7961, 7820, 7681, 7546, 7413,
7282, 7154, 7029, 6906, 6784, 6666, 6551, 6439, 6328, 6219, 6113, 6008, 5906, 5807, 5709, 5613,
5519, 5427, 5337, 5249, 5163, 5079, 4996, 4915, 4836, 4759, 4683, 4608, 4535, 4464, 4394, 4326,
4259, 4193, 4129, 4066, 4004, 3944, 3885, 3827, 3769, 3714, 3660, 3606, 3554, 3502, 3452, 3402,
3354, 3306, 3259, 3214, 3169, 3125, 3082, 3040, 2999, 2958, 2918, 2879, 2840, 2803, 2766, 2729,
2693, 2658, 2624, 2590, 2557, 2525, 2493, 2461, 2430, 2400, 2370, 2341, 2312, 2284, 2256, 2229),
(16266, 16261, 16246, 16220, 16185, 16141, 16086, 16023, 15950, 15867, 15777, 15678, 15570, 15457, 15334, 15206,
15071, 14929, 14782, 14630, 14473, 14310, 14145, 13976, 13803, 13628, 13450, 13270, 13088, 12905, 12720, 12534,
12350, 12164, 11978, 11792, 11607, 11423, 11240, 11057, 10877, 10697, 10519, 10343, 10169, 9997, 9827, 9659,
9493, 9329, 9168, 9009, 8853, 8699, 8547, 8398, 8252, 8108, 7967, 7828, 7691, 7557, 7426, 7296,
7170, 7045, 6925, 6805, 6687, 6574, 6461, 6351, 6243, 6137, 6034, 5932, 5833, 5735, 5640, 5546,
5455, 5365, 5277, 5191, 5107, 5024, 4943, 4864, 4787, 4711, 4636, 4563, 4492, 4422, 4353, 4286,
4220, 4156, 4093, 4031, 3970, 3911, 3853, 3796, 3740, 3685, 3631, 3578, 3527, 3476, 3426, 3377,
3330, 3283, 3237, 3191, 3148, 3105, 3062, 3020, 2979, 2939, 2900, 2861, 2823, 2786, 2749, 2713,
2678, 2643, 2609, 2576, 2543, 2511, 2479, 2448, 2418, 2388, 2358, 2329, 2301, 2273, 2245, 2218),
(15709, 15705, 15691, 15667, 15634, 15593, 15542, 15483, 15415, 15337, 15253, 15161, 15061, 14954, 14840, 14718,
14592, 14460, 14321, 14179, 14030, 13879, 13722, 13564, 13400, 13235, 13067, 12897, 12726, 12552, 12378, 12202,
12026, 11850, 11674, 11497, 11321, 11146, 10971, 10798, 10625, 10454, 10284, 10116, 9949, 9784, 9621, 9460,
9301, 9144, 8989, 8836, 8685, 8537, 8391, 8248, 8105, 7967, 7831, 7697, 7564, 7435, 7308, 7183,
7060, 6940, 6822, 6705, 6592, 6481, 6372, 6265, 6159, 6056, 5956, 5857, 5760, 5665, 5571, 5480,
5391, 5303, 5217, 5133, 5051, 4970, 4891, 4813, 4737, 4663, 4590, 4518, 4448, 4380, 4313, 4247,
4182, 4119, 4057, 3996, 3936, 3878, 3821, 3765, 3710, 3656, 3603, 3551, 3500, 3450, 3401, 3352,
3306, 3259, 3215, 3170, 3127, 3084, 3042, 3001, 2960, 2921, 2882, 2843, 2806, 2769, 2733, 2697,
2663, 2628, 2595, 2562, 2529, 2497, 2466, 2435, 2405, 2375, 2346, 2317, 2289, 2262, 2234, 2208),
(15182, 15176, 15164, 15142, 15112, 15073, 15025, 14970, 14906, 14834, 14754, 14668, 14574, 14474, 14368, 14255,
14136, 14011, 13882, 13747, 13608, 13465, 13318, 13168, 13014, 12859, 12700, 12539, 12377, 12213, 12048, 11881,
11714, 11547, 11379, 11212, 11044, 10877, 10711, 10546, 10381, 10217, 10055, 9894, 9734, 9576, 9420, 9266,
9113, 8962, 8813, 8666, 8522, 8379, 8238, 8100, 7963, 7829, 7697, 7568, 7439, 7315, 7191, 7070,
6952, 6834, 6720, 6608, 6498, 6389, 6283, 6179, 6077, 5976, 5878, 5782, 5687, 5594, 5504, 5415,
5327, 5242, 5158, 5075, 4995, 4916, 4838, 4763, 4688, 4615, 4544, 4474, 4405, 4338, 4272, 4207,
4144, 4082, 4021, 3961, 3902, 3845, 3789, 3733, 3679, 3626, 3574, 3522, 3472, 3424, 3376, 3327,
3282, 3237, 3191, 3148, 3105, 3063, 3021, 2981, 2941, 2902, 2863, 2826, 2789, 2752, 2716, 2681,
2647, 2613, 2580, 2547, 2515, 2484, 2453, 2422, 2392, 2363, 2334, 2306, 2278, 2250, 2223, 2197),
(14680, 14676, 14663, 14643, 14614, 14578, 14534, 14481, 14421, 14355, 14281, 14199, 14112, 14018, 13916, 13811,
13700, 13583, 13461, 13333, 13203, 13069, 12931, 12789, 12644, 12497, 12347, 12195, 12041, 11886, 11729, 11572,
11413, 11254, 11095, 10936, 10776, 10617, 10459, 10301, 10144, 9988, 9832, 9678, 9526, 9374, 9225, 9076,
8930, 8785, 8642, 8500, 8361, 8224, 8087, 7955, 7822, 7693, 7566, 7441, 7317, 7196, 7077, 6959,
6844, 6730, 6619, 6511, 6404, 6299, 6195, 6094, 5995, 5897, 5801, 5707, 5615, 5525, 5436, 5349,
5264, 5180, 5098, 5018, 4939, 4862, 4786, 4712, 4639, 4568, 4498, 4429, 4362, 4296, 4231, 4168,
4105, 4043, 3984, 3926, 3868, 3812, 3757, 3701, 3649, 3597, 3546, 3495, 3445, 3398, 3350, 3304,
3258, 3213, 3169, 3126, 3084, 3042, 3001, 2961, 2922, 2883, 2845, 2808, 2771, 2735, 2700, 2665,
2631, 2598, 2565, 2533, 2501, 2470, 2439, 2409, 2379, 2350, 2322, 2294, 2266, 2239, 2212, 2186),
(14202, 14199, 14187, 14168, 14141, 14107, 14065, 14016, 13961, 13898, 13827, 13752, 13669, 13582, 13488, 13388,
13283, 13173, 13058, 12939, 12816, 12689, 12559, 12425, 12289, 12149, 12008, 11864, 11718, 11571, 11423, 11273,
11123, 10972, 10820, 10669, 10517, 10365, 10214, 10064, 9914, 9764, 9616, 9469, 9322, 9177, 9034, 8892,
8751, 8612, 8474, 8338, 8204, 8072, 7940, 7811, 7685, 7560, 7437, 7316, 7197, 7079, 6963, 6850,
6739, 6629, 6521, 6415, 6311, 6209, 6109, 6010, 5913, 5818, 5725, 5634, 5544, 5456, 5369, 5285,
5201, 5120, 5040, 4961, 4884, 4809, 4734, 4662, 4590, 4520, 4452, 4385, 4319, 4254, 4190, 4128,
4067, 4007, 3948, 3891, 3834, 3778, 3725, 3671, 3619, 3567, 3517, 3468, 3419, 3370, 3325, 3279,
3234, 3190, 3146, 3104, 3062, 3021, 2981, 2941, 2902, 2864, 2827, 2790, 2754, 2718, 2683, 2649,
2615, 2582, 2550, 2518, 2487, 2456, 2426, 2396, 2367, 2338, 2310, 2282, 2254, 2228, 2201, 2175),
(13748, 13744, 13733, 13716, 13691, 13658, 13619, 13574, 13521, 13463, 13397, 13325, 13249, 13166, 13077, 12983,
12885, 12781, 12673, 12561, 12445, 12325, 12202, 12076, 11947, 11815, 11681, 11545, 11407, 11268, 11127, 10985,
10842, 10698, 10554, 10410, 10266, 10121, 9977, 9833, 9690, 9547, 9405, 9264, 9124, 8985, 8848, 8711,
8576, 8442, 8310, 8179, 8050, 7922, 7797, 7673, 7550, 7430, 7310, 7194, 7078, 6965, 6852, 6743,
6635, 6528, 6424, 6321, 6220, 6121, 6023, 5927, 5833, 5741, 5650, 5561, 5473, 5387, 5303, 5220,
5139, 5059, 4981, 4904, 4829, 4755, 4683, 4612, 4542, 4473, 4406, 4340, 4276, 4212, 4150, 4089,
4029, 3970, 3913, 3855, 3800, 3746, 3692, 3640, 3589, 3538, 3488, 3440, 3392, 3345, 3299, 3254,
3209, 3166, 3123, 3081, 3040, 3000, 2960, 2921, 2883, 2845, 2808, 2772, 2736, 2701, 2667, 2633,
2600, 2567, 2535, 2503, 2472, 2442, 2412, 2383, 2354, 2325, 2297, 2270, 2243, 2216, 2190, 2164),
(13314, 13311, 13300, 13285, 13261, 13231, 13195, 13152, 13102, 13047, 12986, 12919, 12845, 12767, 12684, 12597,
12504, 12406, 12304, 12199, 12089, 11976, 11860, 11741, 11619, 11494, 11367, 11238, 11107, 10975, 10842, 10707,
10571, 10434, 10297, 10160, 10022, 9885, 9747, 9610, 9473, 9336, 9201, 9066, 8932, 8798, 8666, 8535,
8406, 8277, 8150, 8024, 7900, 7777, 7656, 7536, 7418, 7301, 7187, 7073, 6962, 6852, 6744, 6637,
6532, 6429, 6328, 6228, 6130, 6033, 5939, 5845, 5754, 5664, 5575, 5489, 5403, 5320, 5237, 5157,
5077, 5000, 4923, 4848, 4775, 4702, 4631, 4562, 4494, 4427, 4361, 4296, 4233, 4171, 4110, 4050,
3991, 3932, 3877, 3821, 3767, 3713, 3660, 3608, 3558, 3509, 3460, 3411, 3365, 3318, 3274, 3229,
3185, 3143, 3100, 3059, 3019, 2979, 2939, 2901, 2863, 2826, 2790, 2754, 2719, 2684, 2650, 2617,
2584, 2552, 2520, 2489, 2458, 2428, 2398, 2369, 2341, 2312, 2285, 2258, 2231, 2205, 2179, 2153),
(12902, 12899, 12889, 12874, 12852, 12823, 12789, 12749, 12702, 12650, 12592, 12530, 12461, 12388, 12309, 12226,
12139, 12047, 11951, 11851, 11748, 11641, 11531, 11418, 11303, 11185, 11065, 10943, 10819, 10693, 10566, 10438,
10309, 10179, 10049, 9918, 9787, 9655, 9524, 9393, 9262, 9132, 9002, 8872, 8744, 8616, 8490, 8364,
8239, 8116, 7993, 7872, 7753, 7634, 7517, 7402, 7288, 7176, 7065, 6955, 6847, 6741, 6636, 6533,
6431, 6331, 6233, 6136, 6041, 5947, 5855, 5764, 5675, 5588, 5502, 5417, 5334, 5252, 5172, 5094,
5016, 4940, 4866, 4792, 4720, 4650, 4581, 4512, 4446, 4380, 4316, 4252, 4190, 4129, 4068, 4011,
3953, 3896, 3841, 3786, 3733, 3680, 3629, 3578, 3528, 3479, 3431, 3384, 3338, 3293, 3248, 3204,
3161, 3119, 3078, 3037, 2997, 2957, 2919, 2881, 2844, 2807, 2771, 2736, 2701, 2667, 2633, 2600,
2568, 2536, 2505, 2474, 2444, 2414, 2385, 2356, 2328, 2300, 2272, 2245, 2219, 2193, 2167, 2142),
(12508, 12505, 12496, 12481, 12461, 12434, 12402, 12364, 12320, 12271, 12217, 12158, 12093, 12024, 11950, 11872,
11789, 11703, 11612, 11518, 11420, 11319, 11216, 11109, 10999, 10888, 10774, 10658, 10540, 10421, 10301, 10179,
10056, 9932, 9808, 9683, 9558, 9433, 9308, 9182, 9057, 8932, 8808, 8684, 8561, 8439, 8317, 8196,
8076, 7958, 7840, 7724, 7609, 7495, 7382, 7271, 7160, 7052, 6945, 6839, 6734, 6632, 6530, 6430,
6332, 6235, 6140, 6046, 5953, 5862, 5772, 5684, 5598, 5513, 5429, 5346, 5266, 5186, 5108, 5031,
4956, 4881, 4809, 4737, 4667, 4598, 4530, 4463, 4398, 4334, 4271, 4209, 4148, 4088, 4029, 3972,
3914, 3860, 3805, 3752, 3699, 3648, 3597, 3547, 3497, 3450, 3403, 3357, 3311, 3266, 3223, 3179,
3137, 3095, 3055, 3014, 2975, 2936, 2898, 2861, 2824, 2788, 2752, 2718, 2683, 2650, 2616, 2584,
2552, 2520, 2489, 2459, 2429, 2400, 2371, 2342, 2314, 2287, 2260, 2233, 2207, 2181, 2156, 2131),
(12132, 12129, 12121, 12107, 12087, 12062, 12032, 11996, 11955, 11909, 11858, 11802, 11742, 11676, 11607, 11533,
11455, 11373, 11287, 11198, 11106, 11010, 10912, 10811, 10707, 10602, 10494, 10384, 10272, 10159, 10044, 9928,
9811, 9694, 9575, 9456, 9337, 9217, 9098, 8978, 8858, 8739, 8620, 8501, 8383, 8266, 8149, 8033,
7918, 7804, 7691, 7579, 7468, 7358, 7249, 7142, 7036, 6931, 6827, 6725, 6623, 6524, 6426, 6329,
6234, 6140, 6047, 5956, 5866, 5778, 5691, 5605, 5521, 5438, 5357, 5277, 5198, 5120, 5044, 4969,
4895, 4823, 4752, 4682, 4613, 4546, 4480, 4414, 4350, 4288, 4226, 4165, 4106, 4047, 3990, 3932,
3878, 3823, 3769, 3717, 3666, 3615, 3565, 3515, 3468, 3420, 3374, 3329, 3284, 3240, 3197, 3155,
3113, 3072, 3032, 2992, 2953, 2915, 2878, 2841, 2804, 2769, 2734, 2699, 2666, 2632, 2600, 2567,
2536, 2505, 2474, 2444, 2415, 2385, 2357, 2329, 2301, 2274, 2247, 2221, 2195, 2170, 2144, 2120),
(11773, 11770, 11762, 11749, 11731, 11707, 11678, 11645, 11606, 11563, 11515, 11462, 11405, 11343, 11277, 11207,
11134, 11056, 10976, 10891, 10804, 10714, 10620, 10525, 10427, 10326, 10224, 10119, 10013, 9905, 9796, 9686,
9575, 9463, 9350, 9237, 9123, 9008, 8894, 8780, 8665, 8551, 8437, 8323, 8210, 8097, 7985, 7874,
7763, 7654, 7545, 7437, 7330, 7224, 7119, 7016, 6913, 6812, 6712, 6612, 6515, 6419, 6324, 6230,
6138, 6047, 5957, 5868, 5781, 5695, 5611, 5527, 5445, 5365, 5285, 5207, 5131, 5055, 4981, 4908,
4836, 4765, 4696, 4627, 4560, 4494, 4430, 4366, 4303, 4242, 4181, 4122, 4064, 4006, 3950, 3895,
3839, 3787, 3734, 3683, 3632, 3581, 3533, 3485, 3438, 3392, 3345, 3300, 3257, 3214, 3171, 3130,
3089, 3048, 3009, 2970, 2931, 2894, 2857, 2820, 2785, 2750, 2715, 2681, 2648, 2615, 2583, 2551,
2520, 2489, 2459, 2429, 2400, 2371, 2343, 2315, 2288, 2261, 2235, 2209, 2183, 2158, 2133, 2109),
(11429, 11426, 11419, 11407, 11389, 11367, 11340, 11308, 11272, 11231, 11185, 11136, 11082, 11024, 10961, 10895,
10826, 10753, 10676, 10597, 10514, 10428, 10340, 10249, 10156, 10061, 9963, 9864, 9763, 9661, 9557, 9452,
9346, 9240, 9132, 9024, 8915, 8806, 8696, 8587, 8477, 8368, 8259, 8150, 8040, 7933, 7826, 7718,
7613, 7507, 7402, 7298, 7195, 7093, 6992, 6891, 6793, 6696, 6598, 6503, 6408, 6315, 6223, 6133,
6043, 5955, 5868, 5782, 5697, 5614, 5531, 5450, 5371, 5292, 5215, 5139, 5064, 4991, 4918, 4847,
4777, 4708, 4640, 4573, 4508, 4443, 4380, 4318, 4257, 4196, 4137, 4079, 4022, 3966, 3910, 3855,
3803, 3750, 3699, 3648, 3599, 3549, 3502, 3454, 3408, 3361, 3318, 3274, 3230, 3188, 3146, 3105,
3064, 3025, 2986, 2947, 2910, 2873, 2836, 2800, 2765, 2730, 2696, 2663, 2630, 2598, 2566, 2534,
2504, 2473, 2443, 2414, 2385, 2357, 2329, 2302, 2275, 2248, 2222, 2196, 2171, 2146, 2121, 2097),
(11100, 11098, 11091, 11079, 11063, 11042, 11016, 10986, 10952, 10913, 10870, 10823, 10772, 10717, 10659, 10596,
10530, 10461, 10389, 10313, 10235, 10154, 10070, 9984, 9895, 9805, 9712, 9618, 9522, 9425, 9326, 9226,
9125, 9023, 8921, 8817, 8714, 8609, 8505, 8400, 8295, 8190, 8086, 7981, 7877, 7772, 7670, 7567,
7464, 7364, 7263, 7163, 7063, 6965, 6868, 6771, 6676, 6580, 6487, 6395, 6304, 6214, 6125, 6037,
5950, 5864, 5780, 5696, 5614, 5533, 5453, 5375, 5297, 5221, 5145, 5071, 4999, 4927, 4856, 4787,
4718, 4651, 4585, 4520, 4456, 4393, 4331, 4270, 4210, 4151, 4093, 4036, 3980, 3925, 3871, 3818,
3766, 3714, 3664, 3614, 3565, 3517, 3470, 3424, 3377, 3333, 3289, 3246, 3204, 3162, 3121, 3080,
3040, 3001, 2963, 2925, 2888, 2851, 2815, 2780, 2745, 2711, 2678, 2645, 2612, 2580, 2549, 2518,
2487, 2458, 2428, 2399, 2371, 2343, 2315, 2288, 2261, 2235, 2209, 2184, 2159, 2134, 2110, 2086),
(10785, 10783, 10776, 10765, 10750, 10730, 10706, 10678, 10645, 10609, 10568, 10524, 10475, 10423, 10368, 10309,
10247, 10181, 10112, 10041, 9967, 9890, 9810, 9728, 9644, 9558, 9471, 9381, 9290, 9197, 9103, 9008,
8911, 8814, 8716, 8618, 8518, 8419, 8319, 8218, 8118, 8018, 7917, 7817, 7717, 7618, 7518, 7420,
7321, 7224, 7127, 7030, 6934, 6840, 6746, 6653, 6561, 6469, 6379, 6290, 6201, 6114, 6028, 5942,
5858, 5775, 5693, 5612, 5532, 5454, 5376, 5300, 5224, 5150, 5077, 5005, 4934, 4864, 4795, 4727,
4661, 4595, 4530, 4467, 4404, 4343, 4282, 4223, 4164, 4106, 4050, 3994, 3939, 3885, 3832, 3780,
3728, 3678, 3629, 3580, 3531, 3485, 3438, 3393, 3348, 3304, 3261, 3219, 3177, 3136, 3095, 3055,
3016, 2978, 2940, 2903, 2866, 2830, 2795, 2760, 2726, 2692, 2659, 2626, 2594, 2563, 2532, 2501,
2471, 2442, 2413, 2384, 2356, 2328, 2301, 2274, 2248, 2222, 2196, 2171, 2146, 2122, 2098, 2075),
(10483, 10481, 10475, 10465, 10450, 10431, 10409, 10382, 10351, 10317, 10278, 10236, 10191, 10141, 10089, 10033,
9974, 9912, 9847, 9779, 9708, 9635, 9560, 9482, 9403, 9321, 9237, 9152, 9065, 8977, 8887, 8796,
8704, 8612, 8518, 8424, 8329, 8234, 8137, 8042, 7946, 7850, 7754, 7657, 7562, 7466, 7371, 7276,
7181, 7087, 6994, 6901, 6809, 6716, 6627, 6537, 6448, 6360, 6272, 6186, 6100, 6016, 5932, 5850,
5768, 5687, 5608, 5529, 5452, 5375, 5300, 5226, 5152, 5080, 5009, 4939, 4870, 4802, 4734, 4668,
4603, 4539, 4476, 4414, 4353, 4293, 4234, 4176, 4118, 4062, 4006, 3952, 3898, 3845, 3793, 3742,
3692, 3642, 3594, 3546, 3499, 3453, 3408, 3363, 3318, 3275, 3232, 3191, 3150, 3110, 3070, 3031,
2992, 2954, 2917, 2880, 2844, 2809, 2774, 2740, 2706, 2673, 2640, 2608, 2576, 2545, 2515, 2485,
2455, 2426, 2397, 2369, 2341, 2314, 2287, 2261, 2235, 2209, 2184, 2159, 2134, 2110, 2086, 2063),
(10194, 10192, 10186, 10177, 10163, 10145, 10124, 10098, 10069, 10036, 10000, 9960, 9917, 9871, 9821, 9768,
9712, 9653, 9591, 9527, 9460, 9391, 9319, 9245, 9169, 9091, 9012, 8931, 8848, 8764, 8678, 8592,
8504, 8416, 8326, 8236, 8144, 8054, 7963, 7871, 7779, 7686, 7593, 7502, 7410, 7317, 7226, 7135,
7044, 6954, 6864, 6773, 6686, 6597, 6510, 6422, 6337, 6252, 6168, 6084, 6001, 5919, 5838, 5758,
5679, 5601, 5524, 5448, 5373, 5298, 5225, 5153, 5082, 5011, 4942, 4874, 4806, 4740, 4675, 4610,
4547, 4484, 4423, 4362, 4302, 4244, 4186, 4129, 4073, 4018, 3963, 3910, 3857, 3805, 3755, 3705,
3656, 3607, 3558, 3513, 3466, 3420, 3376, 3333, 3289, 3247, 3205, 3164, 3123, 3084, 3044, 3006,
2968, 2931, 2894, 2858, 2823, 2788, 2753, 2720, 2686, 2654, 2621, 2590, 2559, 2528, 2498, 2468,
2439, 2410, 2382, 2354, 2327, 2300, 2273, 2247, 2221, 2196, 2171, 2146, 2122, 2098, 2075, 2052),
(9917, 9915, 9909, 9900, 9887, 9870, 9850, 9826, 9798, 9768, 9733, 9695, 9654, 9610, 9563, 9513,
9460, 9404, 9345, 9284, 9221, 9155, 9087, 9016, 8944, 8870, 8794, 8717, 8638, 8558, 8477, 8394,
8310, 8226, 8140, 8054, 7967, 7879, 7792, 7704, 7616, 7528, 7439, 7351, 7262, 7174, 7086, 6998,
6911, 6823, 6737, 6651, 6565, 6480, 6396, 6312, 6229, 6146, 6065, 5984, 5904, 5825, 5746, 5669,
5592, 5516, 5442, 5368, 5295, 5222, 5151, 5081, 5012, 4943, 4876, 4809, 4744, 4679, 4615, 4553,
4491, 4430, 4370, 4310, 4252, 4195, 4138, 4083, 4028, 3973, 3921, 3869, 3817, 3766, 3717, 3667,
3619, 3572, 3524, 3479, 3434, 3389, 3345, 3302, 3259, 3218, 3177, 3137, 3097, 3058, 3019, 2981,
2944, 2907, 2871, 2836, 2801, 2767, 2733, 2699, 2667, 2634, 2603, 2572, 2541, 2511, 2481, 2452,
2423, 2394, 2366, 2339, 2312, 2285, 2259, 2233, 2208, 2183, 2158, 2134, 2110, 2086, 2063, 2040),
(9651, 9649, 9644, 9635, 9622, 9607, 9587, 9565, 9539, 9509, 9477, 9441, 9402, 9360, 9315, 9268,
9217, 9164, 9108, 9050, 8990, 8927, 8863, 8796, 8727, 8657, 8584, 8511, 8436, 8359, 8281, 8202,
8122, 8042, 7960, 7878, 7795, 7711, 7627, 7543, 7457, 7373, 7288, 7203, 7119, 7034, 6949, 6865,
6780, 6697, 6612, 6530, 6447, 6365, 6283, 6203, 6123, 6043, 5964, 5886, 5809, 5732, 5656, 5581,
5507, 5433, 5360, 5289, 5218, 5148, 5078, 5010, 4943, 4876, 4811, 4746, 4682, 4619, 4557, 4496,
4435, 4376, 4317, 4259, 4202, 4146, 4091, 4037, 3982, 3930, 3878, 3827, 3777, 3726, 3679, 3631,
3583, 3537, 3490, 3445, 3401, 3358, 3315, 3272, 3231, 3190, 3148, 3110, 3070, 3032, 2994, 2957,
2920, 2884, 2849, 2814, 2779, 2745, 2712, 2679, 2647, 2615, 2584, 2553, 2523, 2493, 2464, 2435,
2406, 2378, 2351, 2324, 2297, 2271, 2245, 2219, 2194, 2169, 2145, 2121, 2097, 2074, 2051, 2029),
(9395, 9393, 9388, 9380, 9368, 9353, 9335, 9313, 9289, 9261, 9230, 9196, 9159, 9119, 9077, 9032,
8984, 8933, 8880, 8825, 8768, 8708, 8646, 8583, 8518, 8450, 8382, 8311, 8240, 8167, 8092, 8017,
7940, 7863, 7785, 7706, 7627, 7546, 7467, 7385, 7305, 7223, 7142, 7060, 6977, 6897, 6815, 6734,
6653, 6572, 6492, 6412, 6332, 6253, 6175, 6096, 6019, 5942, 5866, 5790, 5715, 5641, 5567, 5494,
5422, 5351, 5281, 5211, 5142, 5074, 5007, 4940, 4875, 4810, 4746, 4683, 4621, 4560, 4499, 4439,
4380, 4322, 4265, 4209, 4153, 4098, 4045, 3991, 3939, 3887, 3837, 3786, 3737, 3689, 3641, 3594,
3547, 3502, 3456, 3413, 3369, 3326, 3284, 3241, 3200, 3161, 3122, 3083, 3044, 3006, 2969, 2932,
2896, 2861, 2826, 2792, 2758, 2724, 2692, 2659, 2627, 2596, 2565, 2535, 2505, 2476, 2447, 2418,
2390, 2363, 2335, 2309, 2282, 2256, 2231, 2205, 2181, 2156, 2132, 2108, 2085, 2062, 2038, 2017),
(9149, 9148, 9143, 9135, 9124, 9110, 9092, 9072, 9049, 9022, 8993, 8961, 8926, 8888, 8847, 8804,
8759, 8711, 8661, 8608, 8553, 8497, 8438, 8377, 8315, 8251, 8186, 8118, 8050, 7980, 7908, 7836,
7764, 7691, 7616, 7539, 7464, 7388, 7310, 7233, 7155, 7077, 6999, 6920, 6841, 6764, 6685, 6607,
6529, 6451, 6374, 6297, 6220, 6143, 6067, 5992, 5917, 5843, 5769, 5696, 5623, 5551, 5480, 5409,
5340, 5271, 5202, 5135, 5068, 5002, 4936, 4872, 4808, 4745, 4683, 4621, 4561, 4501, 4442, 4384,
4326, 4270, 4214, 4159, 4105, 4050, 3998, 3946, 3895, 3845, 3794, 3746, 3698, 3649, 3603, 3556,
3512, 3467, 3422, 3379, 3336, 3295, 3253, 3213, 3172, 3132, 3094, 3056, 3018, 2981, 2944, 2908,
2873, 2838, 2803, 2769, 2736, 2703, 2671, 2639, 2608, 2577, 2547, 2517, 2487, 2458, 2430, 2402,
2374, 2347, 2320, 2293, 2267, 2242, 2217, 2192, 2167, 2143, 2119, 2096, 2073, 2050, 2028, 2006),
(8913, 8912, 8907, 8900, 8889, 8876, 8859, 8840, 8818, 8792, 8765, 8734, 8701, 8665, 8626, 8586,
8542, 8497, 8449, 8399, 8347, 8293, 8237, 8179, 8119, 8058, 7996, 7932, 7867, 7800, 7732, 7664,
7593, 7523, 7452, 7378, 7306, 7233, 7159, 7085, 7010, 6934, 6859, 6784, 6709, 6634, 6558, 6483,
6408, 6333, 6258, 6184, 6110, 6036, 5963, 5890, 5817, 5746, 5674, 5603, 5533, 5463, 5394, 5326,
5258, 5191, 5125, 5059, 4994, 4930, 4867, 4804, 4742, 4681, 4620, 4560, 4501, 4443, 4386, 4329,
4273, 4218, 4163, 4109, 4056, 4004, 3953, 3902, 3852, 3802, 3753, 3706, 3658, 3612, 3565, 3521,
3476, 3433, 3389, 3347, 3305, 3264, 3223, 3182, 3144, 3105, 3066, 3029, 2992, 2955, 2919, 2884,
2849, 2815, 2781, 2747, 2715, 2682, 2651, 2619, 2588, 2558, 2528, 2499, 2470, 2441, 2413, 2385,
2358, 2331, 2304, 2278, 2253, 2227, 2202, 2178, 2154, 2130, 2106, 2083, 2060, 2037, 2016, 1994),
(8686, 8685, 8681, 8673, 8663, 8650, 8635, 8616, 8595, 8571, 8545, 8516, 8484, 8450, 8414, 8375,
8333, 8290, 8244, 8197, 8147, 8096, 8043, 7987, 7931, 7872, 7813, 7752, 7689, 7625, 7561, 7495,
7428, 7360, 7292, 7223, 7153, 7083, 7012, 6940, 6869, 6797, 6725, 6652, 6580, 6507, 6435, 6362,
6290, 6218, 6145, 6074, 6002, 5931, 5860, 5790, 5720, 5650, 5581, 5513, 5445, 5377, 5310, 5244,
5178, 5113, 5049, 4985, 4922, 4860, 4798, 4737, 4677, 4617, 4558, 4500, 4443, 4386, 4330, 4275,
4220, 4166, 4113, 4059, 4009, 3957, 3907, 3858, 3809, 3760, 3713, 3666, 3620, 3574, 3529, 3485,
3441, 3398, 3356, 3314, 3273, 3232, 3193, 3154, 3115, 3077, 3039, 3002, 2966, 2930, 2894, 2860,
2825, 2792, 2758, 2725, 2693, 2661, 2630, 2599, 2569, 2539, 2509, 2480, 2452, 2424, 2396, 2369,
2342, 2315, 2289, 2263, 2238, 2213, 2188, 2164, 2140, 2117, 2093, 2071, 2048, 2026, 2003, 1982),
(8468, 8466, 8462, 8455, 8446, 8434, 8419, 8401, 8381, 8359, 8333, 8306, 8276, 8243, 8208, 8171,
8132, 8091, 8047, 8001, 7955, 7906, 7854, 7802, 7747, 7693, 7636, 7577, 7518, 7457, 7395, 7332,
7267, 7203, 7138, 7070, 7004, 6937, 6869, 6800, 6730, 6662, 6593, 6523, 6454, 6383, 6314, 6244,
6174, 6105, 6035, 5966, 5897, 5828, 5760, 5692, 5624, 5557, 5490, 5424, 5358, 5293, 5228, 5164,
5100, 5037, 4974, 4913, 4851, 4791, 4731, 4671, 4613, 4555, 4497, 4441, 4385, 4329, 4275, 4221,
4168, 4115, 4063, 4012, 3961, 3912, 3862, 3814, 3766, 3719, 3672, 3626, 3581, 3537, 3493, 3449,
3407, 3364, 3323, 3282, 3241, 3202, 3163, 3124, 3086, 3049, 3012, 2976, 2940, 2905, 2870, 2836,
2802, 2769, 2736, 2704, 2672, 2641, 2610, 2579, 2549, 2520, 2491, 2462, 2434, 2406, 2379, 2352,
2325, 2299, 2274, 2248, 2223, 2198, 2174, 2150, 2127, 2103, 2080, 2058, 2036, 2014, 1992, 1970),
(8257, 8256, 8252, 8246, 8237, 8225, 8211, 8194, 8175, 8154, 8130, 8103, 8075, 8044, 8011, 7975,
7938, 7899, 7857, 7814, 7768, 7722, 7673, 7623, 7572, 7519, 7464, 7407, 7351, 7292, 7234, 7174,
7112, 7049, 6988, 6924, 6859, 6795, 6730, 6664, 6598, 6531, 6465, 6397, 6331, 6263, 6196, 6129,
6062, 5995, 5928, 5861, 5794, 5728, 5662, 5596, 5531, 5466, 5401, 5337, 5273, 5210, 5147, 5085,
5023, 4962, 4901, 4841, 4782, 4723, 4664, 4607, 4550, 4493, 4437, 4382, 4328, 4274, 4221, 4168,
4116, 4065, 4014, 3964, 3914, 3866, 3818, 3771, 3724, 3678, 3632, 3587, 3543, 3499, 3456, 3413,
3372, 3331, 3290, 3250, 3209, 3171, 3132, 3095, 3058, 3021, 2985, 2949, 2914, 2879, 2845, 2812,
2778, 2746, 2713, 2682, 2651, 2620, 2589, 2559, 2530, 2501, 2472, 2444, 2416, 2389, 2362, 2335,
2309, 2283, 2258, 2233, 2208, 2184, 2160, 2136, 2113, 2090, 2068, 2045, 2023, 2002, 1980, 1959),
(8055, 8054, 8050, 8044, 8035, 8024, 8011, 7994, 7976, 7956, 7933, 7908, 7881, 7851, 7820, 7786,
7750, 7713, 7673, 7632, 7589, 7545, 7498, 7450, 7401, 7350, 7298, 7245, 7190, 7135, 7078, 7020,
6962, 6902, 6841, 6780, 6719, 6657, 6594, 6531, 6468, 6404, 6340, 6275, 6211, 6146, 6081, 6017,
5952, 5887, 5823, 5758, 5694, 5630, 5566, 5502, 5439, 5376, 5314, 5251, 5190, 5128, 5068, 5007,
4947, 4888, 4829, 4771, 4713, 4656, 4599, 4543, 4487, 4432, 4378, 4324, 4271, 4219, 4167, 4116,
4065, 4015, 3966, 3917, 3869, 3821, 3774, 3728, 3682, 3637, 3592, 3549, 3505, 3462, 3420, 3379,
3338, 3297, 3257, 3218, 3179, 3141, 3103, 3066, 3030, 2994, 2958, 2923, 2888, 2854, 2821, 2788,
2755, 2723, 2691, 2660, 2629, 2599, 2569, 2540, 2511, 2482, 2454, 2426, 2399, 2372, 2345, 2319,
2293, 2268, 2243, 2218, 2194, 2170, 2146, 2123, 2100, 2077, 2055, 2033, 2011, 1989, 1968, 1948),
(7858, 7858, 7854, 7849, 7840, 7829, 7817, 7802, 7785, 7765, 7743, 7720, 7693, 7666, 7636, 7603,
7570, 7534, 7496, 7457, 7416, 7373, 7328, 7283, 7235, 7187, 7138, 7086, 7034, 6981, 6927, 6870,
6815, 6758, 6700, 6642, 6583, 6523, 6463, 6401, 6340, 6279, 6218, 6156, 6094, 6032, 5969, 5907,
5845, 5782, 5720, 5658, 5595, 5534, 5472, 5410, 5349, 5288, 5228, 5168, 5108, 5049, 4990, 4931,
4873, 4815, 4758, 4701, 4645, 4590, 4535, 4480, 4426, 4373, 4320, 4268, 4216, 4165, 4114, 4064,
4015, 3966, 3918, 3870, 3823, 3777, 3731, 3685, 3641, 3597, 3553, 3510, 3468, 3426, 3385, 3343,
3304, 3264, 3225, 3186, 3148, 3111, 3074, 3038, 3002, 2966, 2931, 2897, 2863, 2829, 2796, 2764,
2732, 2700, 2669, 2638, 2608, 2578, 2549, 2520, 2491, 2463, 2435, 2408, 2381, 2355, 2328, 2303,
2277, 2252, 2227, 2203, 2179, 2155, 2132, 2109, 2086, 2064, 2042, 2020, 1998, 1977, 1956, 1935),
(7671, 7670, 7667, 7661, 7653, 7643, 7631, 7617, 7600, 7582, 7561, 7538, 7513, 7486, 7457, 7427,
7395, 7360, 7325, 7287, 7248, 7206, 7165, 7121, 7076, 7030, 6981, 6933, 6883, 6832, 6780, 6727,
6673, 6619, 6562, 6507, 6450, 6393, 6335, 6277, 6218, 6159, 6100, 6040, 5980, 5920, 5860, 5800,
5740, 5680, 5619, 5559, 5499, 5440, 5380, 5321, 5261, 5203, 5144, 5086, 5028, 4970, 4913, 4856,
4800, 4744, 4688, 4633, 4579, 4525, 4471, 4418, 4366, 4314, 4262, 4211, 4161, 4111, 4062, 4013,
3965, 3917, 3870, 3824, 3778, 3733, 3688, 3644, 3599, 3556, 3513, 3472, 3431, 3390, 3349, 3309,
3270, 3231, 3193, 3155, 3118, 3081, 3045, 3009, 2974, 2939, 2905, 2871, 2837, 2805, 2772, 2740,
2709, 2678, 2647, 2617, 2587, 2558, 2529, 2500, 2472, 2444, 2417, 2390, 2364, 2337, 2312, 2286,
2261, 2236, 2212, 2188, 2164, 2141, 2118, 2095, 2073, 2050, 2029, 2007, 1986, 1965, 1944, 1924),
(7489, 7489, 7485, 7480, 7473, 7463, 7451, 7438, 7421, 7403, 7384, 7363, 7339, 7313, 7285, 7257,
7226, 7192, 7159, 7123, 7086, 7047, 7006, 6963, 6920, 6877, 6831, 6784, 6737, 6687, 6637, 6587,
6535, 6483, 6430, 6376, 6321, 6265, 6211, 6155, 6098, 6042, 5984, 5927, 5869, 5812, 5754, 5696,
5638, 5579, 5521, 5463, 5405, 5348, 5290, 5233, 5175, 5118, 5062, 5005, 4949, 4893, 4838, 4783,
4728, 4674, 4620, 4567, 4514, 4461, 4409, 4357, 4306, 4256, 4206, 4156, 4107, 4058, 4009, 3963,
3916, 3870, 3824, 3778, 3733, 3689, 3645, 3602, 3558, 3517, 3475, 3434, 3394, 3354, 3314, 3275,
3236, 3198, 3161, 3124, 3087, 3051, 3016, 2981, 2946, 2912, 2878, 2845, 2812, 2780, 2748, 2717,
2686, 2655, 2625, 2595, 2566, 2537, 2509, 2481, 2453, 2426, 2399, 2372, 2346, 2320, 2295, 2270,
2245, 2221, 2197, 2173, 2149, 2126, 2104, 2081, 2059, 2037, 2016, 1995, 1974, 1952, 1933, 1913),
(7314, 7313, 7310, 7305, 7298, 7289, 7278, 7265, 7249, 7233, 7214, 7192, 7171, 7146, 7120, 7092,
7063, 7031, 6999, 6963, 6929, 6891, 6852, 6813, 6771, 6729, 6685, 6640, 6594, 6548, 6500, 6451,
6401, 6351, 6300, 6249, 6196, 6143, 6090, 6036, 5982, 5927, 5872, 5817, 5761, 5706, 5650, 5594,
5538, 5482, 5426, 5370, 5314, 5258, 5202, 5147, 5091, 5036, 4981, 4926, 4872, 4818, 4764, 4711,
4658, 4605, 4553, 4501, 4449, 4398, 4348, 4298, 4248, 4199, 4150, 4102, 4054, 4006, 3960, 3913,
3868, 3821, 3777, 3733, 3689, 3646, 3603, 3561, 3519, 3478, 3437, 3397, 3357, 3318, 3279, 3241,
3203, 3166, 3129, 3093, 3057, 3022, 2987, 2953, 2919, 2885, 2852, 2819, 2787, 2755, 2724, 2693,
2663, 2633, 2603, 2574, 2545, 2517, 2489, 2461, 2434, 2407, 2380, 2354, 2329, 2303, 2278, 2253,
2229, 2205, 2181, 2158, 2135, 2112, 2090, 2067, 2046, 2024, 2003, 1982, 1961, 1941, 1921, 1901),
(7145, 7144, 7141, 7137, 7130, 7121, 7111, 7098, 7084, 7067, 7049, 7030, 7008, 6984, 6959, 6933,
6905, 6875, 6844, 6811, 6777, 6741, 6704, 6666, 6626, 6585, 6544, 6501, 6457, 6412, 6365, 6319,
6272, 6223, 6174, 6125, 6074, 6024, 5972, 5920, 5868, 5815, 5763, 5709, 5656, 5602, 5548, 5494,
5440, 5386, 5332, 5278, 5224, 5170, 5116, 5062, 5009, 4955, 4902, 4849, 4796, 4744, 4692, 4640,
4589, 4537, 4487, 4436, 4386, 4337, 4287, 4239, 4190, 4142, 4095, 4048, 4000, 3955, 3910, 3864,
3820, 3776, 3732, 3689, 3646, 3604, 3562, 3520, 3479, 3438, 3399, 3360, 3321, 3283, 3245, 3207,
3170, 3134, 3098, 3062, 3027, 2993, 2958, 2925, 2891, 2858, 2826, 2794, 2762, 2731, 2700, 2670,
2640, 2611, 2581, 2553, 2524, 2496, 2469, 2442, 2415, 2388, 2362, 2337, 2311, 2286, 2261, 2237,
2213, 2189, 2166, 2143, 2120, 2098, 2076, 2054, 2032, 2011, 1990, 1969, 1949, 1929, 1909, 1889),
(6981, 6981, 6977, 6974, 6967, 6959, 6949, 6937, 6923, 6908, 6890, 6872, 6851, 6829, 6805, 6779,
6752, 6723, 6694, 6662, 6630, 6594, 6560, 6523, 6485, 6446, 6406, 6365, 6322, 6279, 6236, 6191,
6146, 6099, 6052, 6004, 5956, 5907, 5858, 5808, 5758, 5707, 5656, 5605, 5553, 5501, 5449, 5397,
5345, 5293, 5241, 5188, 5136, 5084, 5032, 4980, 4928, 4876, 4825, 4773, 4722, 4671, 4621, 4571,
4521, 4471, 4422, 4373, 4324, 4276, 4228, 4181, 4134, 4086, 4041, 3995, 3950, 3905, 3860, 3816,
3773, 3728, 3687, 3645, 3603, 3562, 3521, 3479, 3440, 3401, 3361, 3324, 3286, 3248, 3211, 3173,
3138, 3102, 3067, 3032, 2998, 2964, 2930, 2897, 2864, 2832, 2800, 2769, 2738, 2707, 2677, 2647,
2617, 2588, 2560, 2532, 2504, 2476, 2449, 2422, 2396, 2370, 2344, 2319, 2294, 2269, 2245, 2221,
2197, 2174, 2151, 2128, 2105, 2083, 2062, 2040, 2019, 1998, 1977, 1957, 1936, 1917, 1897, 1878),
(6823, 6823, 6821, 6816, 6809, 6802, 6791, 6780, 6768, 6753, 6737, 6719, 6698, 6678, 6655, 6630,
6605, 6576, 6549, 6519, 6487, 6454, 6421, 6385, 6349, 6312, 6272, 6234, 6193, 6152, 6110, 6067,
6023, 5978, 5933, 5887, 5841, 5794, 5746, 5698, 5650, 5601, 5552, 5502, 5453, 5403, 5353, 5302,
5252, 5202, 5151, 5101, 5050, 5000, 4949, 4899, 4849, 4799, 4749, 4699, 4650, 4600, 4551, 4502,
4454, 4406, 4358, 4310, 4263, 4216, 4170, 4124, 4077, 4032, 3987, 3943, 3898, 3855, 3811, 3769,
3726, 3684, 3642, 3601, 3560, 3520, 3479, 3441, 3402, 3363, 3325, 3287, 3250, 3213, 3177, 3141,
3106, 3071, 3036, 3002, 2968, 2935, 2902, 2869, 2837, 2806, 2774, 2743, 2713, 2683, 2653, 2624,
2595, 2566, 2538, 2511, 2483, 2456, 2429, 2403, 2377, 2351, 2326, 2301, 2276, 2252, 2228, 2205,
2181, 2158, 2135, 2113, 2091, 2069, 2048, 2026, 2004, 1985, 1964, 1944, 1924, 1905, 1884, 1866),
(6672, 6671, 6668, 6664, 6658, 6651, 6641, 6630, 6618, 6604, 6587, 6571, 6551, 6532, 6510, 6486,
6462, 6436, 6408, 6379, 6349, 6318, 6285, 6252, 6217, 6181, 6144, 6106, 6068, 6028, 5987, 5946,
5904, 5861, 5818, 5773, 5729, 5683, 5638, 5592, 5545, 5498, 5451, 5403, 5355, 5307, 5258, 5210,
5161, 5113, 5064, 5015, 4966, 4917, 4869, 4820, 4771, 4723, 4674, 4626, 4578, 4530, 4483, 4436,
4389, 4342, 4295, 4249, 4203, 4158, 4112, 4067, 4023, 3979, 3935, 3891, 3848, 3805, 3762, 3722,
3680, 3639, 3598, 3558, 3518, 3479, 3440, 3401, 3363, 3326, 3288, 3252, 3215, 3179, 3144, 3108,
3074, 3039, 3005, 2972, 2939, 2906, 2874, 2842, 2811, 2779, 2749, 2718, 2689, 2659, 2630, 2601,
2573, 2545, 2517, 2490, 2463, 2436, 2410, 2384, 2358, 2333, 2308, 2284, 2259, 2235, 2212, 2188,
2165, 2143, 2120, 2098, 2076, 2055, 2034, 2012, 1992, 1972, 1951, 1932, 1912, 1893, 1873, 1855),
(6524, 6524, 6521, 6517, 6511, 6504, 6494, 6485, 6473, 6458, 6444, 6428, 6410, 6390, 6369, 6347,
6322, 6297, 6272, 6244, 6216, 6186, 6154, 6122, 6089, 6054, 6019, 5983, 5945, 5907, 5868, 5829,
5788, 5747, 5705, 5663, 5620, 5576, 5532, 5488, 5443, 5397, 5352, 5306, 5260, 5213, 5166, 5120,
5073, 5026, 4978, 4931, 4884, 4837, 4790, 4742, 4695, 4648, 4602, 4555, 4508, 4462, 4416, 4370,
4324, 4279, 4234, 4189, 4144, 4100, 4056, 4012, 3969, 3926, 3883, 3841, 3799, 3757, 3716, 3675,
3635, 3595, 3555, 3515, 3477, 3438, 3400, 3363, 3325, 3289, 3252, 3216, 3181, 3145, 3110, 3076,
3042, 3008, 2975, 2942, 2910, 2878, 2846, 2815, 2784, 2754, 2723, 2694, 2664, 2635, 2607, 2578,
2550, 2523, 2496, 2469, 2442, 2416, 2390, 2365, 2340, 2315, 2290, 2266, 2242, 2219, 2195, 2172,
2150, 2127, 2105, 2083, 2062, 2041, 2020, 1999, 1978, 1958, 1939, 1918, 1900, 1880, 1862, 1842),
(6382, 6381, 6379, 6375, 6369, 6362, 6354, 6344, 6332, 6320, 6304, 6289, 6272, 6253, 6233, 6212,
6189, 6165, 6140, 6114, 6086, 6057, 6027, 5996, 5964, 5931, 5897, 5862, 5827, 5790, 5753, 5715,
5676, 5636, 5596, 5555, 5514, 5472, 5429, 5386, 5343, 5299, 5255, 5211, 5166, 5122, 5077, 5031,
4986, 4940, 4895, 4849, 4804, 4758, 4712, 4667, 4621, 4576, 4530, 4485, 4440, 4395, 4350, 4305,
4261, 4217, 4173, 4129, 4086, 4043, 4000, 3957, 3916, 3873, 3832, 3791, 3750, 3710, 3669, 3630,
3590, 3551, 3512, 3474, 3436, 3398, 3361, 3324, 3288, 3252, 3216, 3181, 3146, 3112, 3078, 3044,
3011, 2978, 2945, 2913, 2881, 2850, 2819, 2788, 2758, 2728, 2698, 2669, 2640, 2612, 2584, 2556,
2528, 2501, 2474, 2448, 2422, 2396, 2371, 2346, 2321, 2297, 2272, 2249, 2225, 2202, 2179, 2156,
2134, 2112, 2090, 2069, 2046, 2026, 2006, 1985, 1965, 1944, 1926, 1906, 1887, 1867, 1850, 1831),
(6244, 6243, 6241, 6237, 6232, 6225, 6217, 6208, 6197, 6184, 6170, 6155, 6139, 6121, 6102, 6081,
6059, 6036, 6012, 5987, 5960, 5933, 5904, 5874, 5844, 5812, 5779, 5746, 5711, 5676, 5640, 5604,
5566, 5528, 5489, 5450, 5410, 5370, 5329, 5288, 5246, 5204, 5161, 5119, 5076, 5032, 4989, 4945,
4901, 4857, 4813, 4769, 4725, 4681, 4637, 4592, 4548, 4504, 4460, 4416, 4373, 4329, 4286, 4242,
4199, 4156, 4114, 4071, 4029, 3987, 3946, 3904, 3862, 3821, 3782, 3742, 3701, 3662, 3623, 3583,
3546, 3508, 3470, 3433, 3395, 3359, 3323, 3287, 3250, 3216, 3181, 3146, 3112, 3079, 3045, 3012,
2980, 2947, 2915, 2884, 2853, 2822, 2791, 2761, 2732, 2702, 2673, 2645, 2616, 2588, 2561, 2533,
2506, 2480, 2453, 2428, 2402, 2377, 2352, 2327, 2302, 2278, 2255, 2231, 2208, 2185, 2163, 2140,
2118, 2097, 2075, 2054, 2033, 2012, 1992, 1972, 1952, 1932, 1913, 1893, 1875, 1856, 1838, 1820),
(6110, 6109, 6107, 6104, 6099, 6092, 6085, 6076, 6065, 6053, 6040, 6025, 6010, 5992, 5974, 5954,
5934, 5911, 5888, 5864, 5839, 5812, 5785, 5756, 5726, 5696, 5665, 5633, 5600, 5566, 5531, 5496,
5460, 5423, 5386, 5348, 5310, 5271, 5231, 5192, 5151, 5111, 5070, 5029, 4987, 4945, 4903, 4861,
4819, 4776, 4734, 4691, 4648, 4605, 4563, 4520, 4477, 4434, 4392, 4349, 4307, 4264, 4222, 4180,
4138, 4097, 4055, 4014, 3973, 3932, 3892, 3852, 3812, 3771, 3733, 3692, 3655, 3615, 3578, 3540,
3503, 3465, 3428, 3392, 3356, 3320, 3284, 3249, 3214, 3180, 3146, 3112, 3079, 3046, 3013, 2981,
2949, 2917, 2886, 2855, 2824, 2794, 2764, 2735, 2706, 2677, 2648, 2620, 2593, 2565, 2538, 2511,
2485, 2458, 2433, 2407, 2382, 2357, 2332, 2308, 2284, 2260, 2237, 2214, 2191, 2169, 2146, 2124,
2103, 2081, 2060, 2038, 2019, 1998, 1978, 1958, 1939, 1918, 1900, 1881, 1863, 1844, 1825, 1807),
(5981, 5980, 5978, 5975, 5970, 5964, 5956, 5948, 5938, 5926, 5914, 5900, 5884, 5868, 5850, 5831,
5811, 5790, 5768, 5745, 5720, 5695, 5668, 5641, 5613, 5584, 5553, 5522, 5491, 5458, 5425, 5391,
5356, 5321, 5285, 5249, 5212, 5174, 5136, 5098, 5059, 5020, 4980, 4941, 4901, 4860, 4820, 4779,
4738, 4697, 4656, 4614, 4573, 4531, 4490, 4449, 4407, 4366, 4324, 4283, 4242, 4201, 4160, 4119,
4079, 4038, 3998, 3957, 3918, 3878, 3839, 3800, 3760, 3722, 3684, 3646, 3608, 3570, 3533, 3496,
3460, 3422, 3386, 3352, 3316, 3281, 3247, 3212, 3178, 3145, 3111, 3078, 3046, 3013, 2981, 2950,
2918, 2887, 2857, 2826, 2797, 2767, 2738, 2709, 2680, 2652, 2624, 2596, 2569, 2542, 2515, 2489,
2463, 2437, 2412, 2387, 2362, 2337, 2313, 2289, 2266, 2242, 2219, 2197, 2174, 2152, 2130, 2108,
2087, 2066, 2045, 2025, 2003, 1984, 1964, 1944, 1926, 1906, 1888, 1868, 1850, 1832, 1815, 1797),
(5856, 5855, 5853, 5850, 5845, 5839, 5832, 5824, 5814, 5803, 5791, 5778, 5763, 5747, 5730, 5712,
5693, 5673, 5652, 5629, 5606, 5581, 5556, 5530, 5502, 5474, 5445, 5416, 5385, 5354, 5322, 5289,
5256, 5222, 5187, 5152, 5116, 5080, 5044, 5007, 4969, 4931, 4893, 4855, 4816, 4777, 4738, 4699,
4659, 4619, 4579, 4539, 4499, 4459, 4419, 4379, 4339, 4299, 4259, 4219, 4179, 4139, 4099, 4059,
4020, 3981, 3941, 3903, 3864, 3825, 3787, 3749, 3710, 3673, 3636, 3599, 3562, 3524, 3488, 3453,
3417, 3382, 3347, 3311, 3277, 3243, 3209, 3175, 3143, 3110, 3077, 3045, 3013, 2981, 2950, 2919,
2888, 2858, 2828, 2798, 2769, 2740, 2711, 2683, 2655, 2627, 2599, 2572, 2546, 2519, 2493, 2467,
2441, 2416, 2391, 2367, 2342, 2318, 2294, 2271, 2248, 2225, 2202, 2180, 2157, 2136, 2114, 2093,
2072, 2051, 2029, 2010, 1990, 1969, 1951, 1931, 1912, 1893, 1875, 1857, 1838, 1821, 1803, 1785),
(5734, 5734, 5732, 5729, 5724, 5719, 5712, 5704, 5694, 5684, 5672, 5660, 5646, 5630, 5614, 5597,
5578, 5559, 5538, 5517, 5494, 5471, 5446, 5421, 5395, 5368, 5340, 5312, 5282, 5252, 5221, 5190,
5158, 5125, 5092, 5058, 5024, 4989, 4953, 4918, 4882, 4845, 4808, 4771, 4734, 4696, 4658, 4620,
4582, 4543, 4505, 4466, 4427, 4388, 4350, 4311, 4272, 4233, 4194, 4155, 4116, 4077, 4039, 4000,
3962, 3923, 3886, 3848, 3811, 3773, 3735, 3699, 3662, 3624, 3589, 3553, 3517, 3481, 3445, 3411,
3376, 3341, 3307, 3273, 3239, 3206, 3173, 3139, 3107, 3075, 3043, 3012, 2980, 2949, 2919, 2888,
2858, 2829, 2799, 2770, 2741, 2713, 2685, 2657, 2629, 2602, 2575, 2549, 2522, 2496, 2471, 2445,
2420, 2395, 2371, 2346, 2322, 2299, 2275, 2252, 2229, 2207, 2185, 2163, 2141, 2119, 2098, 2077,
2056, 2036, 2016, 1995, 1976, 1956, 1936, 1918, 1899, 1881, 1862, 1844, 1825, 1808, 1790, 1773),
(5617, 5616, 5614, 5611, 5607, 5602, 5595, 5587, 5578, 5568, 5557, 5545, 5531, 5517, 5501, 5485,
5467, 5448, 5429, 5408, 5386, 5364, 5340, 5316, 5291, 5265, 5238, 5210, 5182, 5153, 5124, 5093,
5062, 5031, 4999, 4966, 4933, 4899, 4865, 4831, 4796, 4761, 4725, 4689, 4653, 4617, 4580, 4543,
4506, 4469, 4432, 4394, 4357, 4319, 4282, 4244, 4206, 4168, 4131, 4093, 4055, 4018, 3980, 3943,
3905, 3869, 3832, 3794, 3758, 3722, 3685, 3649, 3614, 3578, 3542, 3506, 3472, 3437, 3403, 3369,
3334, 3300, 3266, 3234, 3200, 3169, 3136, 3104, 3072, 3041, 3010, 2979, 2948, 2918, 2888, 2858,
2829, 2800, 2771, 2742, 2714, 2686, 2659, 2631, 2604, 2578, 2551, 2525, 2499, 2474, 2449, 2424,
2399, 2374, 2350, 2327, 2303, 2280, 2257, 2234, 2211, 2189, 2167, 2146, 2124, 2103, 2082, 2061,
2041, 2020, 2001, 1981, 1961, 1942, 1923, 1905, 1885, 1867, 1850, 1832, 1814, 1797, 1780, 1763),
(5503, 5502, 5500, 5497, 5493, 5488, 5482, 5475, 5466, 5456, 5446, 5434, 5421, 5407, 5392, 5376,
5359, 5341, 5322, 5302, 5281, 5260, 5237, 5214, 5189, 5164, 5139, 5112, 5085, 5057, 5029, 4999,
4970, 4939, 4908, 4877, 4845, 4812, 4780, 4746, 4713, 4679, 4644, 4610, 4575, 4540, 4504, 4469,
4433, 4397, 4361, 4324, 4288, 4252, 4215, 4178, 4142, 4105, 4068, 4032, 3996, 3959, 3923, 3887,
3850, 3814, 3778, 3743, 3707, 3671, 3636, 3601, 3565, 3531, 3497, 3462, 3428, 3394, 3361, 3327,
3293, 3261, 3228, 3196, 3164, 3132, 3100, 3069, 3038, 3007, 2977, 2946, 2917, 2887, 2857, 2828,
2800, 2771, 2743, 2715, 2687, 2660, 2633, 2606, 2580, 2553, 2527, 2502, 2476, 2451, 2427, 2402,
2378, 2354, 2330, 2307, 2284, 2261, 2238, 2216, 2194, 2172, 2150, 2129, 2108, 2087, 2066, 2046,
2026, 2006, 1986, 1967, 1948, 1929, 1910, 1891, 1873, 1855, 1837, 1820, 1802, 1785, 1768, 1751),
(5392, 5391, 5390, 5387, 5383, 5378, 5372, 5365, 5357, 5348, 5337, 5326, 5313, 5300, 5286, 5270,
5254, 5237, 5218, 5199, 5179, 5158, 5137, 5114, 5091, 5067, 5042, 5017, 4990, 4963, 4936, 4908,
4879, 4850, 4820, 4790, 4759, 4728, 4696, 4664, 4631, 4598, 4565, 4532, 4498, 4464, 4430, 4395,
4361, 4326, 4291, 4256, 4220, 4185, 4150, 4114, 4079, 4043, 4007, 3972, 3937, 3902, 3866, 3830,
3796, 3760, 3726, 3691, 3656, 3622, 3587, 3553, 3519, 3485, 3452, 3418, 3385, 3352, 3318, 3286,
3254, 3222, 3190, 3157, 3127, 3096, 3065, 3034, 3004, 2974, 2944, 2914, 2885, 2856, 2827, 2799,
2771, 2743, 2715, 2688, 2661, 2634, 2607, 2581, 2555, 2529, 2504, 2479, 2454, 2429, 2405, 2381,
2357, 2333, 2310, 2287, 2264, 2242, 2219, 2197, 2176, 2154, 2133, 2112, 2091, 2071, 2050, 2029,
2011, 1991, 1972, 1952, 1934, 1915, 1896, 1878, 1859, 1842, 1824, 1807, 1790, 1773, 1756, 1739),
(5285, 5284, 5283, 5280, 5276, 5271, 5266, 5259, 5251, 5242, 5232, 5221, 5209, 5196, 5183, 5168,
5152, 5135, 5118, 5099, 5080, 5060, 5039, 5018, 4995, 4972, 4948, 4924, 4898, 4872, 4846, 4819,
4791, 4763, 4734, 4705, 4675, 4645, 4614, 4583, 4552, 4520, 4488, 4456, 4423, 4390, 4357, 4324,
4290, 4256, 4223, 4189, 4154, 4120, 4086, 4052, 4016, 3982, 3948, 3914, 3880, 3845, 3811, 3777,
3742, 3708, 3674, 3640, 3607, 3573, 3540, 3506, 3472, 3440, 3407, 3375, 3342, 3309, 3277, 3246,
3215, 3182, 3152, 3121, 3091, 3060, 3030, 3000, 2970, 2941, 2912, 2883, 2854, 2826, 2798, 2770,
2742, 2715, 2688, 2661, 2634, 2608, 2582, 2556, 2531, 2505, 2481, 2456, 2431, 2407, 2383, 2360,
2336, 2313, 2290, 2268, 2245, 2223, 2201, 2179, 2158, 2137, 2116, 2095, 2075, 2055, 2035, 2015,
1995, 1976, 1957, 1938, 1919, 1901, 1883, 1865, 1847, 1830, 1812, 1795, 1778, 1761, 1745, 1728),
(5181, 5180, 5179, 5176, 5172, 5168, 5162, 5156, 5148, 5140, 5130, 5119, 5108, 5096, 5082, 5068,
5053, 5037, 5020, 5002, 4984, 4965, 4945, 4924, 4902, 4880, 4857, 4833, 4809, 4784, 4758, 4732,
4705, 4678, 4650, 4622, 4593, 4564, 4535, 4505, 4474, 4444, 4413, 4382, 4350, 4318, 4286, 4254,
4221, 4189, 4156, 4123, 4090, 4057, 4023, 3990, 3957, 3923, 3889, 3857, 3823, 3790, 3756, 3723,
3690, 3657, 3624, 3590, 3558, 3524, 3493, 3460, 3428, 3395, 3364, 3332, 3300, 3268, 3238, 3207,
3175, 3145, 3115, 3085, 3055, 3025, 2995, 2966, 2937, 2908, 2880, 2852, 2823, 2796, 2768, 2741,
2714, 2687, 2660, 2634, 2608, 2582, 2557, 2532, 2507, 2482, 2457, 2433, 2409, 2385, 2362, 2339,
2316, 2293, 2270, 2248, 2226, 2204, 2183, 2162, 2140, 2120, 2099, 2079, 2059, 2038, 2019, 2000,
1980, 1961, 1943, 1924, 1906, 1887, 1870, 1851, 1833, 1816, 1799, 1782, 1765, 1750, 1733, 1717),
(5080, 5079, 5078, 5075, 5072, 5067, 5062, 5056, 5048, 5040, 5031, 5021, 5010, 4998, 4985, 4971,
4957, 4941, 4925, 4908, 4890, 4872, 4852, 4832, 4811, 4790, 4768, 4745, 4722, 4697, 4673, 4648,
4622, 4596, 4569, 4541, 4514, 4486, 4457, 4428, 4399, 4369, 4339, 4309, 4278, 4248, 4217, 4185,
4154, 4122, 4091, 4059, 4027, 3994, 3962, 3930, 3898, 3864, 3833, 3800, 3768, 3735, 3703, 3671,
3638, 3606, 3574, 3542, 3510, 3478, 3445, 3415, 3383, 3352, 3321, 3290, 3259, 3228, 3198, 3168,
3138, 3108, 3078, 3049, 3019, 2990, 2961, 2933, 2904, 2876, 2848, 2821, 2793, 2766, 2739, 2712,
2686, 2660, 2634, 2608, 2582, 2557, 2532, 2507, 2483, 2458, 2434, 2411, 2387, 2364, 2341, 2318,
2295, 2273, 2251, 2229, 2207, 2186, 2165, 2144, 2123, 2103, 2082, 2062, 2042, 2023, 2003, 1984,
1965, 1947, 1927, 1910, 1892, 1874, 1856, 1839, 1821, 1804, 1787, 1771, 1754, 1738, 1722, 1705),
(4981, 4981, 4979, 4977, 4974, 4970, 4964, 4958, 4951, 4943, 4935, 4925, 4914, 4903, 4890, 4877,
4863, 4848, 4833, 4816, 4799, 4781, 4763, 4743, 4723, 4703, 4681, 4659, 4637, 4613, 4590, 4565,
4540, 4515, 4489, 4463, 4436, 4409, 4381, 4353, 4325, 4296, 4267, 4238, 4209, 4179, 4149, 4119,
4088, 4057, 4027, 3996, 3965, 3932, 3902, 3871, 3839, 3808, 3777, 3744, 3714, 3682, 3651, 3619,
3588, 3556, 3524, 3494, 3463, 3432, 3401, 3370, 3340, 3309, 3279, 3248, 3218, 3188, 3159, 3129,
3100, 3071, 3042, 3013, 2984, 2956, 2928, 2900, 2872, 2845, 2817, 2790, 2763, 2737, 2710, 2684,
2658, 2632, 2607, 2582, 2557, 2532, 2507, 2483, 2459, 2435, 2412, 2388, 2365, 2342, 2320, 2297,
2275, 2253, 2231, 2210, 2189, 2167, 2147, 2126, 2106, 2086, 2066, 2046, 2026, 2007, 1987, 1969,
1951, 1932, 1914, 1896, 1878, 1859, 1842, 1825, 1808, 1791, 1774, 1759, 1742, 1726, 1710, 1695),
(4886, 4886, 4884, 4882, 4879, 4875, 4870, 4864, 4857, 4849, 4841, 4832, 4821, 4810, 4799, 4786,
4772, 4758, 4743, 4727, 4711, 4693, 4676, 4657, 4638, 4618, 4597, 4576, 4554, 4532, 4509, 4485,
4461, 4437, 4412, 4386, 4360, 4334, 4307, 4280, 4253, 4225, 4197, 4169, 4140, 4112, 4082, 4052,
4024, 3994, 3964, 3934, 3904, 3873, 3843, 3812, 3783, 3752, 3721, 3691, 3660, 3630, 3599, 3568,
3538, 3506, 3477, 3447, 3416, 3386, 3356, 3326, 3296, 3266, 3237, 3207, 3178, 3148, 3120, 3091,
3063, 3034, 3006, 2978, 2950, 2922, 2895, 2867, 2840, 2813, 2786, 2760, 2734, 2708, 2682, 2656,
2631, 2606, 2581, 2556, 2531, 2507, 2483, 2459, 2436, 2412, 2389, 2366, 2343, 2321, 2299, 2277,
2255, 2233, 2212, 2191, 2170, 2149, 2129, 2108, 2088, 2069, 2049, 2029, 2010, 1991, 1973, 1953,
1935, 1918, 1900, 1882, 1864, 1847, 1830, 1813, 1796, 1779, 1763, 1747, 1731, 1714, 1699, 1684),
(4793, 4793, 4792, 4789, 4786, 4782, 4778, 4772, 4766, 4758, 4750, 4741, 4731, 4721, 4709, 4697,
4684, 4670, 4656, 4641, 4625, 4608, 4591, 4573, 4554, 4535, 4515, 4494, 4473, 4452, 4430, 4407,
4384, 4360, 4336, 4311, 4286, 4261, 4235, 4209, 4183, 4156, 4129, 4101, 4074, 4046, 4018, 3989,
3961, 3932, 3903, 3873, 3845, 3815, 3786, 3756, 3726, 3697, 3667, 3638, 3608, 3578, 3549, 3519,
3488, 3460, 3429, 3400, 3370, 3342, 3311, 3283, 3254, 3225, 3196, 3166, 3139, 3110, 3082, 3054,
3026, 2998, 2971, 2943, 2916, 2889, 2862, 2835, 2809, 2782, 2756, 2730, 2704, 2679, 2654, 2629,
2604, 2579, 2554, 2530, 2506, 2482, 2459, 2435, 2412, 2389, 2367, 2344, 2322, 2300, 2278, 2256,
2235, 2214, 2193, 2172, 2151, 2131, 2111, 2091, 2071, 2052, 2033, 2012, 1995, 1976, 1957, 1939,
1921, 1902, 1884, 1867, 1850, 1833, 1816, 1799, 1782, 1767, 1751, 1735, 1719, 1703, 1688, 1671),
(4703, 4703, 4702, 4700, 4697, 4693, 4688, 4683, 4677, 4670, 4662, 4653, 4644, 4633, 4622, 4610,
4598, 4585, 4571, 4556, 4541, 4525, 4508, 4491, 4473, 4454, 4435, 4415, 4395, 4374, 4353, 4331,
4308, 4285, 4262, 4238, 4214, 4190, 4165, 4140, 4114, 4088, 4062, 4034, 4007, 3981, 3954, 3927,
3898, 3871, 3843, 3815, 3787, 3758, 3730, 3701, 3672, 3642, 3615, 3586, 3556, 3528, 3499, 3470,
3441, 3411, 3384, 3355, 3326, 3298, 3268, 3241, 3212, 3184, 3156, 3128, 3100, 3072, 3045, 3017,
2990, 2963, 2936, 2909, 2882, 2856, 2829, 2803, 2777, 2752, 2726, 2701, 2676, 2651, 2626, 2601,
2577, 2553, 2529, 2505, 2481, 2458, 2435, 2412, 2389, 2367, 2344, 2322, 2301, 2279, 2257, 2236,
2215, 2194, 2174, 2153, 2133, 2113, 2093, 2074, 2054, 2035, 2016, 1997, 1978, 1960, 1942, 1924,
1906, 1889, 1871, 1854, 1837, 1820, 1804, 1787, 1771, 1755, 1739, 1722, 1706, 1692, 1676, 1661),
(4616, 4615, 4614, 4612, 4609, 4606, 4601, 4596, 4590, 4583, 4576, 4567, 4558, 4548, 4538, 4526,
4514, 4502, 4488, 4474, 4459, 4444, 4428, 4411, 4393, 4376, 4357, 4338, 4318, 4298, 4278, 4256,
4235, 4213, 4190, 4167, 4144, 4120, 4096, 4072, 4047, 4022, 3996, 3971, 3945, 3919, 3892, 3864,
3839, 3812, 3784, 3757, 3730, 3701, 3674, 3647, 3619, 3590, 3563, 3535, 3506, 3478, 3450, 3422,
3394, 3366, 3338, 3309, 3282, 3254, 3227, 3198, 3171, 3144, 3116, 3089, 3062, 3035, 3008, 2981,
2954, 2928, 2901, 2875, 2849, 2823, 2798, 2772, 2747, 2721, 2696, 2672, 2647, 2623, 2598, 2574,
2550, 2527, 2503, 2480, 2457, 2434, 2411, 2389, 2366, 2344, 2323, 2301, 2279, 2258, 2237, 2216,
2196, 2175, 2155, 2135, 2115, 2095, 2076, 2057, 2037, 2019, 2000, 1981, 1963, 1944, 1927, 1909,
1892, 1875, 1857, 1840, 1824, 1807, 1790, 1773, 1757, 1742, 1726, 1711, 1695, 1680, 1665, 1650),
(4531, 4530, 4529, 4527, 4525, 4521, 4517, 4512, 4506, 4499, 4492, 4484, 4475, 4466, 4455, 4445,
4433, 4421, 4408, 4394, 4380, 4365, 4349, 4333, 4316, 4299, 4281, 4263, 4244, 4224, 4204, 4184,
4163, 4142, 4120, 4098, 4075, 4052, 4029, 4005, 3981, 3957, 3932, 3907, 3882, 3857, 3830, 3805,
3780, 3753, 3726, 3701, 3674, 3647, 3620, 3592, 3565, 3539, 3512, 3484, 3456, 3429, 3403, 3375,
3348, 3321, 3293, 3266, 3239, 3212, 3185, 3157, 3130, 3104, 3077, 3051, 3024, 2998, 2971, 2945,
2919, 2893, 2868, 2842, 2817, 2791, 2766, 2741, 2716, 2692, 2667, 2643, 2619, 2595, 2571, 2548,
2524, 2501, 2478, 2455, 2433, 2410, 2388, 2366, 2344, 2322, 2301, 2280, 2258, 2238, 2217, 2196,
2176, 2156, 2136, 2116, 2097, 2078, 2058, 2038, 2020, 2002, 1984, 1966, 1948, 1930, 1912, 1895,
1876, 1859, 1842, 1827, 1810, 1794, 1778, 1762, 1746, 1730, 1714, 1699, 1684, 1669, 1654, 1638),
(4448, 4448, 4447, 4445, 4442, 4439, 4435, 4430, 4424, 4418, 4411, 4403, 4394, 4385, 4375, 4365,
4354, 4342, 4329, 4316, 4302, 4288, 4273, 4257, 4241, 4224, 4207, 4189, 4171, 4152, 4133, 4113,
4093, 4072, 4050, 4030, 4007, 3986, 3963, 3939, 3917, 3894, 3870, 3846, 3821, 3796, 3771, 3747,
3722, 3696, 3671, 3645, 3619, 3592, 3567, 3540, 3515, 3488, 3462, 3435, 3409, 3382, 3356, 3329,
3302, 3275, 3249, 3223, 3196, 3170, 3144, 3117, 3091, 3065, 3039, 3013, 2987, 2961, 2936, 2910,
2885, 2859, 2834, 2809, 2784, 2760, 2735, 2711, 2686, 2662, 2638, 2615, 2591, 2568, 2544, 2521,
2498, 2476, 2453, 2431, 2408, 2386, 2365, 2343, 2322, 2300, 2279, 2258, 2238, 2217, 2197, 2177,
2157, 2137, 2118, 2098, 2079, 2060, 2041, 2023, 2003, 1986, 1968, 1950, 1932, 1915, 1897, 1880,
1863, 1846, 1830, 1813, 1797, 1781, 1765, 1748, 1733, 1718, 1702, 1687, 1671, 1657, 1643, 1628),
(4368, 4367, 4366, 4364, 4362, 4358, 4354, 4350, 4344, 4338, 4332, 4324, 4316, 4307, 4297, 4287,
4276, 4265, 4253, 4240, 4227, 4213, 4199, 4184, 4168, 4152, 4135, 4118, 4100, 4082, 4063, 4043,
4025, 4005, 3984, 3964, 3943, 3921, 3898, 3877, 3855, 3832, 3809, 3786, 3762, 3737, 3714, 3690,
3665, 3641, 3615, 3590, 3565, 3540, 3515, 3490, 3463, 3438, 3413, 3386, 3361, 3336, 3309, 3284,
3258, 3232, 3206, 3180, 3155, 3129, 3103, 3078, 3052, 3026, 3001, 2976, 2950, 2925, 2900, 2875,
2851, 2826, 2801, 2777, 2753, 2728, 2704, 2680, 2657, 2633, 2610, 2587, 2563, 2540, 2518, 2495,
2473, 2450, 2428, 2406, 2385, 2363, 2342, 2320, 2299, 2279, 2258, 2237, 2217, 2197, 2177, 2157,
2138, 2118, 2099, 2080, 2061, 2043, 2024, 2006, 1987, 1969, 1952, 1934, 1917, 1900, 1882, 1866,
1849, 1832, 1816, 1799, 1784, 1768, 1752, 1736, 1721, 1705, 1691, 1676, 1661, 1646, 1632, 1617),
(4289, 4289, 4288, 4286, 4284, 4280, 4277, 4272, 4267, 4261, 4254, 4247, 4239, 4231, 4222, 4212,
4201, 4190, 4179, 4166, 4154, 4140, 4126, 4112, 4097, 4081, 4065, 4048, 4031, 4014, 3996, 3977,
3957, 3939, 3919, 3898, 3879, 3858, 3837, 3815, 3794, 3771, 3749, 3726, 3703, 3681, 3657, 3633,
3610, 3586, 3562, 3538, 3513, 3488, 3463, 3440, 3415, 3390, 3365, 3340, 3315, 3290, 3264, 3239,
3214, 3189, 3164, 3139, 3114, 3088, 3063, 3038, 3013, 2989, 2964, 2939, 2915, 2890, 2866, 2841,
2817, 2793, 2769, 2745, 2721, 2698, 2674, 2651, 2628, 2605, 2582, 2559, 2536, 2514, 2491, 2469,
2447, 2426, 2404, 2382, 2361, 2340, 2319, 2298, 2278, 2257, 2237, 2217, 2197, 2177, 2157, 2138,
2119, 2100, 2081, 2062, 2044, 2025, 2007, 1989, 1970, 1953, 1935, 1918, 1901, 1884, 1867, 1850,
1835, 1818, 1802, 1786, 1770, 1755, 1739, 1723, 1709, 1694, 1679, 1663, 1649, 1635, 1620, 1607),
(4213, 4213, 4212, 4210, 4208, 4205, 4201, 4196, 4191, 4186, 4179, 4172, 4165, 4157, 4148, 4138,
4128, 4117, 4106, 4093, 4082, 4068, 4056, 4041, 4027, 4012, 3996, 3980, 3964, 3947, 3929, 3911,
3893, 3875, 3855, 3836, 3816, 3796, 3776, 3755, 3734, 3712, 3691, 3669, 3647, 3624, 3602, 3579,
3556, 3533, 3509, 3486, 3462, 3438, 3413, 3390, 3366, 3342, 3318, 3293, 3268, 3245, 3220, 3196,
3171, 3147, 3122, 3098, 3073, 3049, 3024, 3000, 2976, 2951, 2927, 2903, 2879, 2855, 2831, 2808,
2784, 2760, 2737, 2714, 2690, 2667, 2644, 2621, 2599, 2576, 2554, 2532, 2509, 2487, 2466, 2444,
2422, 2401, 2380, 2359, 2338, 2317, 2297, 2276, 2256, 2236, 2216, 2196, 2177, 2157, 2138, 2119,
2100, 2081, 2063, 2044, 2026, 2008, 1990, 1973, 1955, 1938, 1919, 1902, 1885, 1870, 1853, 1837,
1821, 1804, 1789, 1773, 1756, 1742, 1726, 1711, 1696, 1682, 1667, 1652, 1637, 1624, 1610, 1595),
(4139, 4138, 4137, 4136, 4133, 4131, 4127, 4123, 4118, 4112, 4106, 4100, 4092, 4084, 4075, 4067,
4057, 4047, 4036, 4024, 4012, 4000, 3987, 3973, 3959, 3944, 3929, 3914, 3898, 3880, 3864, 3846,
3830, 3812, 3793, 3774, 3755, 3735, 3716, 3696, 3675, 3655, 3633, 3612, 3590, 3569, 3547, 3524,
3503, 3479, 3458, 3435, 3411, 3389, 3365, 3342, 3318, 3295, 3272, 3248, 3224, 3200, 3177, 3153,
3129, 3105, 3081, 3057, 3033, 3010, 2986, 2962, 2938, 2915, 2891, 2868, 2844, 2821, 2798, 2774,
2751, 2728, 2705, 2683, 2660, 2637, 2615, 2593, 2570, 2548, 2526, 2505, 2483, 2461, 2440, 2419,
2398, 2377, 2356, 2335, 2315, 2294, 2274, 2254, 2234, 2215, 2195, 2176, 2157, 2138, 2119, 2100,
2081, 2063, 2045, 2027, 2009, 1991, 1973, 1956, 1939, 1922, 1905, 1888, 1871, 1855, 1839, 1823,
1807, 1790, 1774, 1760, 1744, 1729, 1714, 1699, 1684, 1670, 1654, 1641, 1627, 1612, 1599, 1585),
(4066, 4066, 4065, 4064, 4061, 4059, 4055, 4050, 4046, 4041, 4034, 4029, 4022, 4014, 4006, 3997,
3987, 3977, 3966, 3956, 3944, 3932, 3920, 3905, 3893, 3879, 3864, 3849, 3834, 3818, 3802, 3785,
3768, 3750, 3732, 3714, 3696, 3676, 3658, 3638, 3617, 3598, 3578, 3556, 3536, 3515, 3494, 3472,
3451, 3429, 3407, 3385, 3363, 3340, 3317, 3295, 3272, 3249, 3225, 3203, 3180, 3157, 3134, 3111,
3087, 3064, 3041, 3018, 2994, 2971, 2948, 2925, 2902, 2879, 2856, 2833, 2810, 2787, 2764, 2742,
2719, 2697, 2674, 2652, 2630, 2608, 2586, 2564, 2542, 2521, 2499, 2478, 2457, 2436, 2415, 2394,
2373, 2353, 2332, 2312, 2292, 2272, 2252, 2233, 2213, 2194, 2175, 2156, 2137, 2118, 2100, 2081,
2063, 2045, 2027, 2009, 1992, 1974, 1957, 1940, 1923, 1906, 1889, 1873, 1856, 1840, 1824, 1807,
1793, 1777, 1762, 1746, 1731, 1716, 1701, 1687, 1671, 1658, 1643, 1629, 1615, 1601, 1587, 1574),
(3996, 3996, 3995, 3993, 3991, 3988, 3984, 3981, 3977, 3972, 3966, 3960, 3953, 3945, 3937, 3929,
3920, 3910, 3900, 3889, 3878, 3866, 3854, 3841, 3828, 3815, 3801, 3786, 3771, 3756, 3740, 3724,
3707, 3690, 3673, 3655, 3637, 3619, 3599, 3581, 3562, 3543, 3522, 3503, 3483, 3463, 3442, 3420,
3400, 3379, 3357, 3336, 3314, 3292, 3270, 3248, 3225, 3204, 3182, 3159, 3137, 3114, 3092, 3069,
3047, 3024, 3001, 2979, 2956, 2933, 2911, 2888, 2866, 2843, 2821, 2798, 2776, 2754, 2732, 2710,
2687, 2666, 2644, 2622, 2600, 2579, 2557, 2536, 2515, 2493, 2472, 2452, 2431, 2410, 2390, 2369,
2349, 2329, 2309, 2289, 2269, 2250, 2231, 2211, 2192, 2173, 2154, 2136, 2117, 2099, 2081, 2063,
2045, 2027, 2009, 1992, 1975, 1957, 1940, 1924, 1907, 1890, 1874, 1858, 1842, 1825, 1810, 1794,
1779, 1763, 1748, 1733, 1718, 1704, 1688, 1674, 1660, 1646, 1632, 1618, 1603, 1590, 1577, 1564),
(3927, 3927, 3926, 3925, 3923, 3920, 3917, 3913, 3909, 3904, 3898, 3892, 3886, 3878, 3871, 3862,
3854, 3844, 3835, 3824, 3812, 3802, 3790, 3778, 3765, 3752, 3737, 3724, 3710, 3694, 3680, 3664,
3648, 3632, 3615, 3598, 3580, 3563, 3545, 3526, 3508, 3488, 3470, 3450, 3431, 3411, 3391, 3370,
3350, 3330, 3309, 3288, 3266, 3246, 3224, 3203, 3181, 3160, 3138, 3116, 3094, 3073, 3051, 3029,
3007, 2985, 2962, 2940, 2918, 2896, 2874, 2852, 2830, 2808, 2786, 2765, 2743, 2721, 2699, 2678,
2656, 2635, 2613, 2592, 2571, 2550, 2529, 2508, 2487, 2467, 2446, 2426, 2405, 2385, 2365, 2345,
2325, 2305, 2286, 2266, 2247, 2228, 2209, 2190, 2171, 2153, 2134, 2116, 2098, 2080, 2062, 2044,
2027, 2009, 1992, 1975, 1958, 1941, 1924, 1908, 1891, 1875, 1859, 1842, 1827, 1811, 1796, 1780,
1765, 1750, 1735, 1720, 1705, 1691, 1677, 1662, 1648, 1634, 1620, 1607, 1593, 1578, 1566, 1553),
(3861, 3860, 3859, 3858, 3855, 3853, 3850, 3846, 3842, 3837, 3832, 3827, 3820, 3812, 3805, 3798,
3789, 3780, 3771, 3760, 3750, 3739, 3728, 3716, 3703, 3691, 3678, 3664, 3649, 3636, 3621, 3606,
3590, 3574, 3558, 3542, 3524, 3508, 3490, 3472, 3454, 3436, 3417, 3399, 3379, 3360, 3341, 3321,
3300, 3281, 3261, 3241, 3221, 3200, 3179, 3157, 3137, 3116, 3095, 3074, 3053, 3031, 3010, 2989,
2967, 2946, 2924, 2903, 2881, 2860, 2838, 2817, 2795, 2774, 2753, 2731, 2710, 2689, 2668, 2647,
2626, 2605, 2584, 2563, 2542, 2522, 2501, 2481, 2460, 2440, 2420, 2400, 2380, 2360, 2341, 2321,
2302, 2282, 2263, 2244, 2225, 2206, 2188, 2169, 2151, 2133, 2114, 2096, 2079, 2061, 2043, 2026,
2009, 1992, 1975, 1958, 1941, 1924, 1908, 1892, 1876, 1859, 1844, 1828, 1812, 1797, 1782, 1765,
1751, 1737, 1722, 1706, 1693, 1678, 1663, 1650, 1636, 1621, 1609, 1595, 1582, 1569, 1555, 1542),
(3794, 3794, 3794, 3793, 3791, 3789, 3786, 3782, 3778, 3773, 3768, 3762, 3756, 3750, 3742, 3735,
3726, 3718, 3709, 3699, 3689, 3678, 3667, 3656, 3644, 3631, 3619, 3605, 3592, 3578, 3564, 3549,
3534, 3519, 3503, 3487, 3470, 3454, 3437, 3420, 3402, 3384, 3366, 3348, 3330, 3311, 3292, 3273,
3254, 3234, 3215, 3195, 3175, 3155, 3135, 3115, 3094, 3074, 3053, 3033, 3012, 2991, 2970, 2949,
2929, 2908, 2887, 2866, 2845, 2824, 2803, 2782, 2761, 2740, 2719, 2699, 2678, 2657, 2636, 2616,
2595, 2575, 2554, 2534, 2514, 2494, 2473, 2454, 2434, 2414, 2394, 2375, 2355, 2336, 2316, 2297,
2278, 2259, 2241, 2222, 2203, 2185, 2167, 2148, 2130, 2112, 2095, 2077, 2060, 2042, 2025, 2008,
1991, 1974, 1957, 1941, 1924, 1908, 1892, 1876, 1859, 1844, 1829, 1813, 1798, 1782, 1768, 1753,
1738, 1722, 1709, 1694, 1680, 1666, 1652, 1637, 1624, 1611, 1597, 1584, 1570, 1558, 1545, 1532),
(3732, 3732, 3731, 3728, 3728, 3725, 3722, 3719, 3715, 3710, 3706, 3700, 3694, 3688, 3681, 3673,
3665, 3657, 3648, 3639, 3629, 3619, 3608, 3597, 3585, 3573, 3561, 3547, 3535, 3521, 3508, 3493,
3479, 3463, 3449, 3433, 3417, 3401, 3385, 3368, 3351, 3334, 3316, 3299, 3281, 3262, 3243, 3225,
3207, 3188, 3169, 3150, 3130, 3111, 3091, 3072, 3052, 3032, 3012, 2992, 2972, 2952, 2931, 2911,
2891, 2870, 2850, 2829, 2809, 2789, 2768, 2748, 2727, 2707, 2687, 2666, 2646, 2626, 2606, 2585,
2565, 2545, 2525, 2506, 2486, 2466, 2446, 2427, 2407, 2388, 2369, 2350, 2330, 2311, 2293, 2274,
2255, 2237, 2218, 2200, 2182, 2164, 2146, 2128, 2110, 2093, 2075, 2058, 2041, 2024, 2007, 1990,
1973, 1957, 1940, 1924, 1908, 1892, 1876, 1859, 1845, 1829, 1814, 1799, 1782, 1769, 1754, 1739,
1723, 1710, 1696, 1682, 1668, 1654, 1640, 1626, 1612, 1599, 1586, 1573, 1560, 1547, 1534, 1521),
(3670, 3670, 3669, 3667, 3666, 3664, 3660, 3657, 3654, 3649, 3644, 3639, 3633, 3626, 3620, 3613,
3605, 3597, 3589, 3580, 3570, 3560, 3549, 3539, 3528, 3515, 3504, 3492, 3479, 3466, 3453, 3438,
3425, 3410, 3395, 3381, 3365, 3350, 3334, 3317, 3300, 3284, 3266, 3250, 3232, 3215, 3197, 3179,
3161, 3143, 3124, 3106, 3087, 3068, 3049, 3030, 3010, 2991, 2972, 2952, 2932, 2913, 2893, 2873,
2853, 2833, 2814, 2794, 2774, 2754, 2734, 2714, 2694, 2674, 2654, 2635, 2615, 2595, 2575, 2556,
2536, 2516, 2497, 2477, 2458, 2439, 2420, 2400, 2381, 2362, 2344, 2325, 2306, 2288, 2269, 2251,
2232, 2214, 2196, 2178, 2160, 2143, 2125, 2108, 2090, 2073, 2056, 2038, 2021, 2004, 1989, 1972,
1956, 1940, 1923, 1907, 1892, 1876, 1859, 1845, 1829, 1814, 1799, 1784, 1769, 1755, 1739, 1725,
1711, 1697, 1683, 1669, 1654, 1641, 1628, 1614, 1601, 1587, 1575, 1562, 1549, 1536, 1524, 1511),
(3610, 3608, 3608, 3607, 3606, 3603, 3601, 3597, 3594, 3590, 3585, 3580, 3574, 3568, 3562, 3555,
3547, 3539, 3531, 3522, 3513, 3503, 3493, 3483, 3472, 3461, 3449, 3437, 3425, 3411, 3399, 3386,
3372, 3358, 3343, 3329, 3314, 3299, 3284, 3268, 3252, 3236, 3219, 3203, 3186, 3169, 3151, 3134,
3116, 3098, 3080, 3062, 3044, 3026, 3007, 2988, 2970, 2951, 2932, 2913, 2894, 2874, 2855, 2836,
2817, 2797, 2778, 2759, 2739, 2720, 2700, 2681, 2661, 2642, 2623, 2603, 2584, 2565, 2545, 2526,
2507, 2488, 2469, 2450, 2431, 2412, 2393, 2374, 2356, 2337, 2319, 2300, 2282, 2264, 2246, 2228,
2210, 2192, 2174, 2157, 2139, 2122, 2105, 2088, 2071, 2054, 2037, 2020, 2003, 1986, 1970, 1955,
1938, 1923, 1907, 1891, 1875, 1859, 1845, 1829, 1814, 1799, 1784, 1770, 1755, 1740, 1726, 1712,
1697, 1684, 1670, 1655, 1643, 1629, 1616, 1603, 1589, 1576, 1563, 1551, 1538, 1525, 1513, 1501),
(3551, 3549, 3549, 3547, 3547, 3545, 3542, 3539, 3535, 3531, 3527, 3522, 3515, 3510, 3504, 3497,
3490, 3483, 3475, 3466, 3456, 3447, 3438, 3428, 3418, 3407, 3395, 3384, 3372, 3360, 3347, 3334,
3321, 3307, 3293, 3279, 3265, 3250, 3234, 3220, 3204, 3188, 3172, 3156, 3139, 3123, 3106, 3089,
3072, 3055, 3037, 3020, 3002, 2984, 2966, 2948, 2930, 2911, 2893, 2874, 2856, 2837, 2818, 2799,
2781, 2762, 2743, 2724, 2705, 2686, 2667, 2648, 2629, 2610, 2591, 2572, 2554, 2535, 2516, 2497,
2478, 2460, 2441, 2422, 2404, 2386, 2367, 2349, 2331, 2312, 2294, 2276, 2258, 2241, 2223, 2205,
2188, 2170, 2153, 2136, 2119, 2101, 2085, 2068, 2051, 2034, 2018, 2002, 1985, 1969, 1952, 1936,
1921, 1906, 1890, 1875, 1859, 1844, 1829, 1814, 1799, 1784, 1770, 1755, 1740, 1727, 1713, 1699,
1685, 1671, 1657, 1644, 1629, 1617, 1603, 1591, 1578, 1565, 1552, 1540, 1527, 1515, 1503, 1490),
(3493, 3493, 3492, 3490, 3488, 3487, 3485, 3481, 3478, 3474, 3470, 3465, 3460, 3454, 3447, 3442,
3435, 3427, 3419, 3411, 3403, 3394, 3384, 3374, 3364, 3354, 3343, 3332, 3320, 3308, 3296, 3283,
3270, 3257, 3243, 3230, 3216, 3202, 3187, 3172, 3157, 3141, 3126, 3111, 3095, 3079, 3062, 3046,
3029, 3012, 2995, 2978, 2961, 2943, 2926, 2908, 2890, 2872, 2854, 2836, 2818, 2800, 2782, 2764,
2745, 2727, 2708, 2690, 2672, 2653, 2635, 2616, 2598, 2579, 2561, 2542, 2524, 2505, 2487, 2469,
2450, 2432, 2414, 2396, 2377, 2359, 2341, 2324, 2306, 2288, 2270, 2253, 2235, 2218, 2200, 2183,
2166, 2149, 2132, 2115, 2098, 2081, 2065, 2048, 2032, 2015, 1999, 1983, 1967, 1951, 1935, 1919,
1904, 1889, 1874, 1859, 1842, 1828, 1814, 1799, 1784, 1770, 1755, 1740, 1727, 1713, 1699, 1685,
1671, 1658, 1645, 1631, 1618, 1604, 1592, 1578, 1566, 1554, 1541, 1529, 1516, 1504, 1492, 1480),
(3437, 3437, 3436, 3435, 3433, 3431, 3429, 3426, 3422, 3419, 3415, 3410, 3404, 3399, 3393, 3386,
3379, 3373, 3366, 3358, 3349, 3341, 3331, 3322, 3311, 3302, 3291, 3281, 3268, 3258, 3246, 3234,
3221, 3207, 3195, 3182, 3168, 3154, 3139, 3126, 3111, 3096, 3081, 3066, 3051, 3035, 3019, 3003,
2987, 2970, 2954, 2937, 2920, 2903, 2886, 2869, 2852, 2834, 2817, 2799, 2782, 2764, 2746, 2728,
2711, 2693, 2675, 2657, 2639, 2621, 2603, 2584, 2566, 2548, 2530, 2512, 2494, 2476, 2458, 2440,
2422, 2405, 2387, 2369, 2351, 2334, 2316, 2299, 2281, 2264, 2246, 2229, 2212, 2195, 2178, 2161,
2144, 2127, 2111, 2094, 2078, 2061, 2045, 2029, 2012, 1997, 1981, 1965, 1949, 1934, 1918, 1902,
1888, 1872, 1857, 1842, 1828, 1813, 1798, 1784, 1770, 1755, 1740, 1727, 1713, 1699, 1686, 1671,
1659, 1645, 1632, 1619, 1606, 1593, 1580, 1568, 1555, 1543, 1530, 1518, 1506, 1494, 1482, 1470),
(3382, 3382, 3381, 3379, 3379, 3377, 3374, 3372, 3368, 3365, 3361, 3356, 3351, 3345, 3340, 3334,
3327, 3320, 3313, 3305, 3297, 3289, 3280, 3271, 3261, 3250, 3241, 3231, 3220, 3207, 3197, 3185,
3173, 3161, 3148, 3135, 3122, 3108, 3094, 3081, 3066, 3052, 3037, 3022, 3007, 2992, 2977, 2961,
2945, 2929, 2913, 2897, 2881, 2864, 2848, 2831, 2814, 2797, 2780, 2763, 2746, 2728, 2711, 2694,
2676, 2659, 2641, 2624, 2606, 2589, 2571, 2553, 2536, 2518, 2501, 2483, 2465, 2448, 2430, 2413,
2395, 2378, 2360, 2343, 2326, 2308, 2291, 2274, 2257, 2240, 2223, 2206, 2189, 2172, 2156, 2139,
2123, 2106, 2090, 2074, 2057, 2041, 2025, 2009, 1994, 1978, 1961, 1947, 1932, 1916, 1901, 1885,
1871, 1856, 1841, 1827, 1812, 1798, 1782, 1769, 1755, 1740, 1727, 1713, 1700, 1686, 1671, 1659,
1646, 1633, 1620, 1607, 1594, 1581, 1569, 1556, 1544, 1531, 1519, 1507, 1495, 1483, 1472, 1460),
(3329, 3329, 3327, 3327, 3325, 3323, 3321, 3318, 3315, 3311, 3308, 3302, 3299, 3293, 3288, 3282,
3275, 3268, 3262, 3254, 3246, 3238, 3230, 3221, 3212, 3202, 3191, 3182, 3171, 3160, 3148, 3138,
3126, 3114, 3102, 3089, 3076, 3063, 3050, 3036, 3022, 3008, 2994, 2980, 2965, 2950, 2935, 2920,
2905, 2889, 2873, 2858, 2842, 2826, 2810, 2793, 2777, 2760, 2744, 2727, 2710, 2694, 2677, 2660,
2643, 2626, 2609, 2591, 2574, 2557, 2540, 2523, 2506, 2488, 2471, 2454, 2437, 2420, 2402, 2385,
2368, 2351, 2334, 2317, 2300, 2283, 2266, 2250, 2233, 2216, 2200, 2183, 2167, 2150, 2134, 2118,
2101, 2085, 2069, 2053, 2037, 2021, 2006, 1990, 1975, 1960, 1944, 1929, 1914, 1899, 1884, 1868,
1854, 1840, 1824, 1811, 1797, 1782, 1768, 1754, 1739, 1727, 1713, 1699, 1686, 1672, 1659, 1646,
1633, 1620, 1607, 1595, 1582, 1569, 1557, 1545, 1532, 1520, 1508, 1496, 1485, 1473, 1461, 1450),
(3277, 3275, 3275, 3275, 3273, 3271, 3268, 3266, 3264, 3259, 3256, 3252, 3247, 3241, 3237, 3231,
3225, 3219, 3212, 3204, 3197, 3189, 3181, 3172, 3163, 3154, 3144, 3134, 3124, 3113, 3102, 3091,
3080, 3068, 3056, 3044, 3031, 3019, 3006, 2993, 2979, 2966, 2952, 2938, 2923, 2909, 2894, 2880,
2865, 2850, 2834, 2819, 2804, 2788, 2772, 2756, 2740, 2724, 2708, 2692, 2676, 2659, 2643, 2626,
2610, 2593, 2576, 2560, 2543, 2526, 2509, 2493, 2476, 2459, 2442, 2425, 2409, 2392, 2375, 2358,
2342, 2325, 2308, 2292, 2275, 2259, 2242, 2226, 2209, 2193, 2177, 2160, 2144, 2128, 2112, 2096,
2080, 2065, 2049, 2033, 2018, 2002, 1986, 1972, 1956, 1941, 1926, 1910, 1897, 1882, 1867, 1853,
1838, 1824, 1810, 1795, 1781, 1767, 1753, 1739, 1726, 1712, 1699, 1686, 1671, 1659, 1646, 1633,
1620, 1608, 1595, 1582, 1569, 1558, 1545, 1533, 1521, 1509, 1498, 1486, 1474, 1463, 1451, 1440),
(3225, 3225, 3225, 3224, 3222, 3221, 3218, 3216, 3213, 3209, 3206, 3202, 3197, 3191, 3187, 3182,
3175, 3169, 3163, 3156, 3148, 3139, 3132, 3124, 3115, 3106, 3097, 3087, 3077, 3067, 3057, 3046,
3035, 3023, 3012, 3000, 2988, 2975, 2963, 2950, 2937, 2924, 2910, 2897, 2883, 2869, 2855, 2840,
2826, 2811, 2796, 2781, 2766, 2751, 2736, 2720, 2705, 2689, 2673, 2657, 2642, 2626, 2610, 2593,
2577, 2561, 2545, 2529, 2512, 2496, 2479, 2463, 2447, 2430, 2414, 2397, 2381, 2365, 2348, 2332,
2315, 2299, 2283, 2267, 2250, 2234, 2218, 2202, 2186, 2170, 2154, 2138, 2122, 2107, 2091, 2075,
2060, 2044, 2029, 2014, 1998, 1983, 1968, 1952, 1938, 1923, 1909, 1893, 1879, 1865, 1850, 1836,
1822, 1807, 1794, 1780, 1765, 1752, 1739, 1725, 1712, 1697, 1685, 1671, 1659, 1646, 1633, 1620,
1608, 1595, 1583, 1569, 1558, 1546, 1534, 1522, 1510, 1498, 1487, 1475, 1464, 1452, 1441, 1430),
(3175, 3175, 3175, 3173, 3173, 3171, 3169, 3166, 3163, 3160, 3157, 3153, 3148, 3144, 3139, 3132,
3127, 3121, 3115, 3108, 3101, 3093, 3085, 3077, 3069, 3060, 3051, 3042, 3032, 3022, 3012, 3001,
2991, 2980, 2968, 2957, 2945, 2933, 2921, 2908, 2896, 2883, 2870, 2856, 2843, 2829, 2816, 2802,
2787, 2773, 2759, 2744, 2729, 2715, 2700, 2685, 2670, 2654, 2639, 2624, 2608, 2592, 2577, 2561,
2545, 2530, 2514, 2498, 2482, 2466, 2450, 2434, 2418, 2402, 2386, 2370, 2354, 2338, 2322, 2306,
2290, 2274, 2258, 2242, 2226, 2210, 2194, 2179, 2163, 2147, 2132, 2116, 2101, 2085, 2070, 2055,
2038, 2024, 2009, 1994, 1978, 1964, 1949, 1935, 1919, 1906, 1891, 1876, 1862, 1848, 1833, 1820,
1806, 1791, 1778, 1765, 1751, 1738, 1723, 1711, 1697, 1685, 1671, 1659, 1646, 1633, 1620, 1608,
1595, 1583, 1570, 1559, 1547, 1535, 1523, 1511, 1499, 1488, 1476, 1465, 1453, 1442, 1431, 1420),
(3127, 3127, 3126, 3125, 3124, 3122, 3120, 3118, 3115, 3112, 3109, 3105, 3100, 3096, 3091, 3086,
3080, 3074, 3068, 3061, 3054, 3047, 3039, 3032, 3023, 3015, 3006, 2997, 2988, 2978, 2968, 2958,
2947, 2937, 2926, 2914, 2903, 2891, 2880, 2867, 2855, 2843, 2830, 2817, 2804, 2791, 2777, 2764,
2750, 2736, 2722, 2708, 2693, 2679, 2664, 2650, 2635, 2620, 2605, 2590, 2575, 2560, 2545, 2529,
2514, 2499, 2483, 2468, 2452, 2436, 2421, 2405, 2390, 2374, 2358, 2343, 2327, 2311, 2296, 2280,
2264, 2249, 2233, 2218, 2202, 2187, 2171, 2156, 2140, 2125, 2110, 2094, 2079, 2064, 2049, 2034,
2019, 2003, 1990, 1975, 1960, 1946, 1931, 1917, 1901, 1888, 1874, 1859, 1846, 1832, 1818, 1804,
1790, 1777, 1763, 1750, 1736, 1722, 1710, 1697, 1684, 1671, 1658, 1645, 1633, 1620, 1608, 1595,
1583, 1570, 1559, 1547, 1535, 1523, 1511, 1500, 1488, 1477, 1465, 1454, 1443, 1432, 1421, 1410),
(3079, 3079, 3079, 3078, 3077, 3075, 3073, 3071, 3068, 3065, 3062, 3058, 3054, 3049, 3045, 3039,
3034, 3028, 3022, 3016, 3009, 3002, 2995, 2987, 2979, 2971, 2962, 2953, 2944, 2935, 2925, 2915,
2905, 2895, 2884, 2873, 2862, 2851, 2839, 2827, 2815, 2803, 2791, 2778, 2766, 2753, 2740, 2726,
2713, 2699, 2686, 2672, 2658, 2644, 2630, 2616, 2601, 2587, 2572, 2558, 2543, 2528, 2513, 2498,
2483, 2468, 2453, 2438, 2423, 2407, 2392, 2377, 2362, 2346, 2331, 2316, 2300, 2285, 2270, 2255,
2239, 2224, 2209, 2194, 2178, 2163, 2148, 2133, 2118, 2103, 2088, 2073, 2058, 2043, 2029, 2014,
1999, 1985, 1969, 1956, 1941, 1927, 1913, 1899, 1884, 1870, 1857, 1842, 1829, 1815, 1801, 1788,
1773, 1761, 1748, 1735, 1721, 1708, 1695, 1683, 1670, 1657, 1644, 1632, 1620, 1607, 1595, 1583,
1570, 1559, 1547, 1535, 1523, 1512, 1500, 1489, 1477, 1466, 1455, 1444, 1433, 1422, 1411, 1400),
(3033, 3033, 3032, 3031, 3030, 3029, 3027, 3024, 3022, 3019, 3016, 3012, 3008, 3004, 2999, 2994,
2989, 2983, 2977, 2971, 2965, 2958, 2951, 2943, 2935, 2927, 2919, 2910, 2902, 2893, 2883, 2874,
2864, 2854, 2843, 2833, 2822, 2811, 2800, 2788, 2776, 2765, 2753, 2740, 2728, 2715, 2703, 2690,
2677, 2664, 2650, 2637, 2623, 2610, 2596, 2582, 2568, 2554, 2540, 2525, 2511, 2497, 2482, 2467,
2453, 2438, 2423, 2409, 2394, 2379, 2364, 2349, 2334, 2319, 2304, 2289, 2274, 2259, 2244, 2230,
2215, 2200, 2185, 2170, 2155, 2140, 2125, 2111, 2096, 2081, 2066, 2052, 2037, 2023, 2008, 1994,
1980, 1965, 1951, 1936, 1923, 1909, 1895, 1881, 1867, 1853, 1840, 1825, 1812, 1799, 1785, 1772,
1759, 1746, 1733, 1720, 1706, 1694, 1680, 1669, 1655, 1644, 1631, 1619, 1607, 1594, 1582, 1569,
1559, 1547, 1535, 1523, 1512, 1500, 1489, 1478, 1467, 1456, 1445, 1434, 1423, 1412, 1401, 1391),
(2988, 2987, 2987, 2986, 2985, 2983, 2981, 2979, 2977, 2974, 2971, 2967, 2963, 2959, 2955, 2950,
2945, 2939, 2934, 2927, 2921, 2914, 2908, 2900, 2893, 2885, 2877, 2869, 2860, 2851, 2842, 2833,
2823, 2813, 2803, 2793, 2782, 2772, 2761, 2750, 2738, 2727, 2715, 2703, 2691, 2679, 2667, 2654,
2641, 2629, 2616, 2603, 2589, 2576, 2563, 2549, 2535, 2522, 2508, 2494, 2480, 2466, 2452, 2437,
2423, 2409, 2394, 2380, 2365, 2351, 2336, 2322, 2307, 2293, 2278, 2263, 2249, 2234, 2220, 2205,
2190, 2176, 2161, 2146, 2132, 2117, 2103, 2088, 2074, 2060, 2045, 2031, 2017, 2002, 1987, 1974,
1960, 1946, 1932, 1918, 1904, 1891, 1876, 1863, 1850, 1836, 1823, 1808, 1796, 1782, 1770, 1756,
1744, 1731, 1718, 1705, 1692, 1680, 1667, 1654, 1642, 1629, 1618, 1606, 1594, 1582, 1569, 1558,
1546, 1535, 1523, 1512, 1500, 1489, 1478, 1467, 1456, 1445, 1434, 1423, 1413, 1402, 1392, 1381),
(2943, 2943, 2942, 2942, 2941, 2939, 2937, 2935, 2933, 2930, 2927, 2923, 2920, 2916, 2911, 2907,
2902, 2896, 2891, 2885, 2879, 2872, 2865, 2858, 2851, 2844, 2836, 2828, 2819, 2811, 2802, 2793,
2783, 2774, 2764, 2754, 2744, 2733, 2723, 2712, 2701, 2690, 2678, 2667, 2655, 2643, 2631, 2619,
2607, 2594, 2582, 2569, 2556, 2543, 2530, 2517, 2503, 2490, 2476, 2463, 2449, 2435, 2422, 2408,
2394, 2380, 2366, 2352, 2338, 2323, 2309, 2295, 2281, 2266, 2252, 2238, 2224, 2209, 2195, 2181,
2166, 2152, 2138, 2123, 2109, 2095, 2081, 2067, 2053, 2037, 2024, 2010, 1995, 1982, 1969, 1955,
1941, 1927, 1913, 1900, 1885, 1873, 1859, 1846, 1833, 1819, 1806, 1793, 1780, 1767, 1754, 1740,
1728, 1716, 1703, 1689, 1678, 1666, 1653, 1641, 1629, 1617, 1604, 1593, 1581, 1569, 1558, 1546,
1534, 1523, 1512, 1500, 1489, 1478, 1467, 1456, 1445, 1434, 1424, 1413, 1403, 1392, 1382, 1372),
(2900, 2900, 2899, 2898, 2897, 2896, 2894, 2892, 2889, 2887, 2884, 2880, 2877, 2873, 2869, 2864,
2859, 2854, 2849, 2843, 2837, 2831, 2824, 2817, 2810, 2803, 2795, 2788, 2779, 2771, 2762, 2754,
2745, 2735, 2726, 2716, 2706, 2696, 2686, 2675, 2664, 2653, 2642, 2631, 2620, 2608, 2596, 2585,
2572, 2560, 2548, 2536, 2523, 2510, 2498, 2485, 2472, 2459, 2446, 2432, 2419, 2406, 2392, 2379,
2365, 2351, 2338, 2324, 2310, 2296, 2282, 2268, 2254, 2241, 2227, 2213, 2199, 2185, 2171, 2157,
2143, 2129, 2115, 2101, 2087, 2073, 2059, 2045, 2031, 2017, 2003, 1990, 1976, 1963, 1949, 1935,
1922, 1908, 1895, 1882, 1867, 1855, 1842, 1829, 1816, 1803, 1790, 1777, 1764, 1751, 1738, 1726,
1713, 1701, 1688, 1676, 1663, 1652, 1638, 1627, 1615, 1603, 1592, 1580, 1568, 1557, 1545, 1534,
1523, 1511, 1500, 1489, 1478, 1467, 1456, 1445, 1435, 1424, 1414, 1403, 1393, 1382, 1372, 1362),
(2857, 2857, 2857, 2856, 2855, 2853, 2852, 2850, 2847, 2845, 2842, 2839, 2835, 2831, 2827, 2823,
2818, 2813, 2808, 2802, 2796, 2790, 2784, 2777, 2770, 2763, 2756, 2748, 2740, 2732, 2724, 2715,
2706, 2697, 2688, 2679, 2669, 2659, 2649, 2639, 2628, 2618, 2607, 2596, 2585, 2574, 2562, 2551,
2539, 2527, 2515, 2503, 2491, 2478, 2466, 2453, 2441, 2428, 2415, 2402, 2389, 2376, 2363, 2350,
2337, 2323, 2310, 2296, 2283, 2269, 2256, 2242, 2229, 2215, 2201, 2188, 2174, 2160, 2147, 2133,
2119, 2106, 2092, 2078, 2065, 2051, 2037, 2024, 2010, 1997, 1983, 1969, 1956, 1943, 1930, 1916,
1902, 1890, 1876, 1864, 1850, 1838, 1824, 1812, 1799, 1786, 1773, 1761, 1748, 1736, 1722, 1711,
1697, 1686, 1674, 1662, 1650, 1637, 1626, 1614, 1602, 1590, 1578, 1567, 1556, 1544, 1533, 1522,
1511, 1500, 1489, 1478, 1467, 1456, 1445, 1435, 1424, 1414, 1403, 1393, 1383, 1373, 1363, 1353),
(2816, 2816, 2815, 2814, 2813, 2812, 2810, 2808, 2806, 2803, 2801, 2798, 2794, 2790, 2786, 2782,
2778, 2773, 2768, 2762, 2757, 2751, 2744, 2738, 2731, 2724, 2717, 2710, 2702, 2694, 2686, 2678,
2669, 2660, 2651, 2642, 2633, 2623, 2613, 2603, 2593, 2583, 2572, 2562, 2551, 2540, 2529, 2518,
2506, 2495, 2483, 2471, 2459, 2447, 2435, 2423, 2410, 2398, 2385, 2373, 2360, 2347, 2335, 2322,
2309, 2296, 2283, 2270, 2256, 2243, 2230, 2217, 2203, 2190, 2177, 2163, 2150, 2137, 2123, 2110,
2096, 2083, 2070, 2056, 2043, 2029, 2016, 2003, 1990, 1976, 1963, 1950, 1936, 1924, 1910, 1898,
1884, 1872, 1859, 1846, 1833, 1820, 1807, 1795, 1782, 1770, 1756, 1745, 1731, 1720, 1708, 1696,
1684, 1671, 1660, 1648, 1636, 1624, 1612, 1601, 1589, 1578, 1566, 1555, 1543, 1532, 1521, 1510,
1499, 1488, 1477, 1467, 1456, 1445, 1435, 1424, 1414, 1404, 1393, 1383, 1373, 1363, 1353, 1343),
(2775, 2775, 2774, 2774, 2773, 2771, 2770, 2768, 2766, 2763, 2760, 2757, 2754, 2750, 2747, 2742,
2738, 2733, 2728, 2723, 2718, 2712, 2706, 2700, 2693, 2686, 2679, 2672, 2665, 2657, 2649, 2641,
2633, 2624, 2615, 2606, 2597, 2588, 2578, 2569, 2559, 2549, 2538, 2528, 2518, 2507, 2496, 2485,
2474, 2463, 2451, 2440, 2428, 2416, 2405, 2393, 2381, 2368, 2356, 2344, 2332, 2319, 2307, 2294,
2281, 2269, 2256, 2243, 2230, 2217, 2204, 2191, 2178, 2165, 2152, 2139, 2126, 2113, 2100, 2087,
2074, 2061, 2048, 2035, 2020, 2008, 1995, 1982, 1969, 1956, 1943, 1930, 1918, 1905, 1892, 1879,
1866, 1854, 1841, 1828, 1816, 1803, 1790, 1778, 1765, 1754, 1740, 1729, 1717, 1705, 1693, 1680,
1669, 1657, 1645, 1634, 1621, 1610, 1599, 1586, 1576, 1565, 1553, 1542, 1531, 1520, 1509, 1498,
1487, 1477, 1466, 1455, 1445, 1434, 1424, 1414, 1404, 1393, 1383, 1373, 1363, 1353, 1344, 1334),
(2735, 2735, 2735, 2734, 2733, 2732, 2730, 2728, 2726, 2724, 2721, 2718, 2715, 2711, 2708, 2704,
2699, 2695, 2690, 2685, 2679, 2674, 2668, 2662, 2656, 2649, 2642, 2635, 2628, 2620, 2613, 2605,
2597, 2588, 2580, 2571, 2562, 2553, 2544, 2534, 2525, 2515, 2505, 2495, 2485, 2474, 2464, 2453,
2442, 2431, 2420, 2409, 2398, 2386, 2375, 2363, 2351, 2339, 2327, 2315, 2303, 2291, 2279, 2267,
2254, 2242, 2229, 2217, 2204, 2192, 2179, 2166, 2154, 2141, 2128, 2116, 2103, 2090, 2077, 2064,
2051, 2038, 2026, 2012, 2000, 1986, 1975, 1961, 1949, 1935, 1924, 1910, 1898, 1885, 1873, 1861,
1848, 1836, 1823, 1811, 1799, 1786, 1773, 1762, 1750, 1738, 1726, 1714, 1702, 1689, 1678, 1666,
1654, 1643, 1631, 1620, 1608, 1597, 1586, 1574, 1563, 1552, 1541, 1530, 1519, 1508, 1497, 1487,
1476, 1465, 1455, 1444, 1434, 1424, 1414, 1403, 1393, 1383, 1373, 1363, 1354, 1344, 1334, 1325),
(2696, 2696, 2696, 2695, 2694, 2693, 2691, 2690, 2687, 2685, 2683, 2680, 2676, 2673, 2669, 2665,
2661, 2657, 2652, 2647, 2642, 2637, 2631, 2625, 2619, 2612, 2606, 2599, 2592, 2585, 2577, 2570,
2562, 2554, 2545, 2537, 2528, 2519, 2510, 2501, 2492, 2482, 2472, 2463, 2453, 2442, 2432, 2422,
2411, 2400, 2390, 2379, 2368, 2356, 2345, 2334, 2322, 2311, 2299, 2288, 2276, 2264, 2252, 2240,
2228, 2216, 2204, 2191, 2179, 2167, 2154, 2142, 2130, 2117, 2105, 2092, 2080, 2067, 2055, 2042,
2029, 2017, 2003, 1992, 1978, 1967, 1953, 1942, 1929, 1917, 1904, 1892, 1880, 1867, 1855, 1842,
1830, 1818, 1806, 1794, 1782, 1770, 1757, 1746, 1734, 1722, 1710, 1697, 1686, 1675, 1663, 1652,
1640, 1629, 1617, 1606, 1595, 1584, 1572, 1561, 1550, 1539, 1528, 1518, 1507, 1496, 1486, 1475,
1465, 1454, 1444, 1433, 1423, 1413, 1403, 1393, 1383, 1373, 1363, 1354, 1344, 1334, 1325, 1315),
(2658, 2658, 2658, 2657, 2656, 2655, 2653, 2652, 2650, 2647, 2645, 2642, 2639, 2636, 2632, 2628,
2624, 2620, 2615, 2610, 2605, 2600, 2595, 2589, 2583, 2577, 2570, 2564, 2557, 2550, 2542, 2535,
2527, 2519, 2511, 2503, 2495, 2486, 2477, 2468, 2459, 2450, 2440, 2431, 2421, 2411, 2401, 2391,
2381, 2370, 2360, 2349, 2338, 2327, 2316, 2305, 2294, 2283, 2271, 2260, 2249, 2237, 2225, 2214,
2202, 2190, 2178, 2166, 2154, 2142, 2130, 2118, 2106, 2094, 2081, 2069, 2057, 2045, 2032, 2020,
2008, 1995, 1983, 1970, 1959, 1946, 1934, 1922, 1910, 1898, 1884, 1873, 1861, 1849, 1837, 1824,
1813, 1801, 1789, 1777, 1765, 1753, 1740, 1730, 1718, 1705, 1695, 1683, 1671, 1660, 1649, 1637,
1626, 1615, 1603, 1592, 1581, 1569, 1559, 1548, 1538, 1527, 1516, 1505, 1495, 1484, 1474, 1464,
1453, 1443, 1433, 1423, 1413, 1403, 1393, 1383, 1373, 1363, 1354, 1344, 1334, 1325, 1316, 1306),
(2621, 2621, 2620, 2620, 2619, 2618, 2616, 2614, 2613, 2610, 2608, 2605, 2602, 2599, 2595, 2592,
2588, 2584, 2579, 2574, 2570, 2564, 2559, 2553, 2548, 2542, 2535, 2529, 2522, 2515, 2508, 2501,
2493, 2486, 2478, 2470, 2462, 2453, 2445, 2436, 2427, 2418, 2409, 2399, 2390, 2380, 2371, 2361,
2351, 2340, 2330, 2320, 2309, 2299, 2288, 2277, 2266, 2255, 2244, 2233, 2222, 2210, 2199, 2188,
2176, 2165, 2153, 2141, 2130, 2118, 2106, 2094, 2082, 2070, 2058, 2046, 2035, 2023, 2011, 1999,
1986, 1974, 1961, 1950, 1938, 1926, 1914, 1901, 1890, 1878, 1866, 1855, 1842, 1831, 1819, 1807,
1795, 1784, 1772, 1760, 1748, 1737, 1725, 1714, 1702, 1691, 1679, 1668, 1657, 1645, 1634, 1623,
1612, 1601, 1590, 1578, 1568, 1557, 1546, 1536, 1525, 1514, 1504, 1493, 1483, 1473, 1462, 1452,
1442, 1432, 1422, 1412, 1402, 1392, 1382, 1373, 1363, 1353, 1344, 1334, 1325, 1316, 1306, 1297),
(2584, 2584, 2584, 2583, 2582, 2581, 2580, 2578, 2576, 2574, 2572, 2569, 2566, 2563, 2560, 2556,
2552, 2548, 2544, 2539, 2534, 2529, 2524, 2519, 2513, 2507, 2501, 2495, 2488, 2482, 2475, 2468,
2460, 2453, 2445, 2437, 2429, 2421, 2413, 2404, 2396, 2387, 2378, 2369, 2360, 2350, 2341, 2331,
2321, 2311, 2301, 2291, 2281, 2271, 2260, 2250, 2239, 2228, 2217, 2206, 2195, 2184, 2173, 2162,
2151, 2140, 2128, 2117, 2105, 2094, 2082, 2071, 2059, 2046, 2036, 2024, 2012, 2001, 1989, 1977,
1965, 1953, 1942, 1930, 1918, 1907, 1895, 1883, 1871, 1859, 1848, 1836, 1824, 1813, 1801, 1790,
1778, 1767, 1755, 1744, 1731, 1721, 1709, 1697, 1687, 1675, 1663, 1653, 1642, 1631, 1620, 1609,
1598, 1586, 1576, 1566, 1555, 1544, 1534, 1523, 1513, 1502, 1492, 1482, 1471, 1461, 1451, 1441,
1431, 1421, 1411, 1401, 1391, 1382, 1372, 1363, 1353, 1344, 1334, 1325, 1316, 1306, 1297, 1288),
(2549, 2548, 2548, 2547, 2547, 2545, 2544, 2543, 2541, 2539, 2536, 2534, 2531, 2528, 2525, 2521,
2517, 2513, 2509, 2505, 2500, 2495, 2490, 2485, 2479, 2474, 2468, 2462, 2455, 2449, 2442, 2435,
2428, 2421, 2413, 2406, 2398, 2390, 2382, 2373, 2365, 2356, 2348, 2339, 2330, 2321, 2311, 2302,
2292, 2283, 2273, 2263, 2253, 2243, 2233, 2222, 2212, 2202, 2191, 2180, 2170, 2159, 2148, 2137,
2126, 2115, 2104, 2093, 2082, 2070, 2059, 2048, 2036, 2025, 2014, 2002, 1991, 1978, 1968, 1956,
1944, 1933, 1922, 1910, 1899, 1887, 1876, 1864, 1851, 1841, 1830, 1818, 1807, 1795, 1784, 1772,
1761, 1750, 1738, 1727, 1716, 1705, 1694, 1682, 1671, 1660, 1649, 1637, 1627, 1617, 1606, 1595,
1584, 1574, 1563, 1552, 1542, 1531, 1521, 1511, 1500, 1490, 1480, 1470, 1460, 1450, 1440, 1430,
1420, 1410, 1400, 1391, 1381, 1371, 1362, 1353, 1343, 1334, 1325, 1315, 1306, 1297, 1288, 1279),
(2514, 2513, 2513, 2512, 2512, 2511, 2509, 2508, 2506, 2504, 2502, 2499, 2496, 2493, 2490, 2487,
2483, 2479, 2475, 2471, 2466, 2462, 2457, 2451, 2446, 2441, 2435, 2429, 2423, 2416, 2410, 2403,
2396, 2389, 2382, 2374, 2367, 2359, 2351, 2343, 2335, 2326, 2318, 2309, 2300, 2291, 2282, 2273,
2264, 2255, 2245, 2235, 2226, 2216, 2206, 2196, 2186, 2175, 2165, 2155, 2144, 2134, 2123, 2112,
2102, 2091, 2080, 2069, 2058, 2046, 2036, 2025, 2014, 2003, 1992, 1980, 1969, 1958, 1947, 1935,
1924, 1913, 1901, 1890, 1879, 1867, 1856, 1845, 1833, 1823, 1811, 1799, 1789, 1778, 1767, 1755,
1744, 1733, 1722, 1711, 1700, 1688, 1678, 1667, 1655, 1645, 1635, 1624, 1612, 1602, 1592, 1581,
1570, 1560, 1550, 1539, 1529, 1519, 1508, 1498, 1488, 1478, 1468, 1458, 1448, 1438, 1428, 1419,
1409, 1399, 1390, 1380, 1371, 1361, 1352, 1343, 1333, 1324, 1315, 1306, 1297, 1288, 1279, 1270),
(2479, 2479, 2479, 2478, 2477, 2476, 2475, 2474, 2472, 2470, 2468, 2465, 2462, 2460, 2456, 2453,
2450, 2446, 2442, 2438, 2433, 2429, 2424, 2419, 2414, 2408, 2403, 2397, 2391, 2385, 2378, 2372,
2365, 2358, 2351, 2344, 2336, 2329, 2321, 2313, 2305, 2297, 2289, 2280, 2272, 2263, 2254, 2245,
2236, 2227, 2218, 2208, 2199, 2189, 2179, 2169, 2160, 2150, 2140, 2129, 2119, 2109, 2098, 2088,
2078, 2067, 2056, 2046, 2035, 2024, 2014, 2003, 1992, 1981, 1969, 1959, 1948, 1936, 1926, 1915,
1904, 1893, 1882, 1871, 1859, 1849, 1838, 1827, 1816, 1805, 1794, 1782, 1771, 1761, 1750, 1739,
1728, 1717, 1705, 1695, 1684, 1672, 1663, 1652, 1641, 1631, 1620, 1609, 1599, 1587, 1578, 1568,
1557, 1547, 1537, 1526, 1516, 1506, 1496, 1486, 1476, 1466, 1456, 1446, 1437, 1427, 1417, 1408,
1398, 1389, 1379, 1370, 1360, 1351, 1342, 1333, 1324, 1315, 1306, 1297, 1288, 1279, 1270, 1262),
(2446, 2445, 2445, 2445, 2444, 2443, 2442, 2440, 2438, 2436, 2434, 2432, 2429, 2427, 2423, 2420,
2417, 2413, 2409, 2405, 2401, 2396, 2392, 2387, 2382, 2376, 2371, 2365, 2359, 2353, 2347, 2341,
2334, 2328, 2321, 2314, 2306, 2299, 2292, 2284, 2276, 2268, 2260, 2252, 2243, 2235, 2226, 2218,
2209, 2200, 2191, 2181, 2172, 2163, 2153, 2144, 2134, 2124, 2114, 2105, 2095, 2084, 2074, 2064,
2054, 2044, 2033, 2023, 2012, 2002, 1991, 1981, 1969, 1959, 1949, 1938, 1927, 1917, 1906, 1895,
1884, 1873, 1863, 1851, 1841, 1830, 1819, 1807, 1797, 1787, 1776, 1765, 1754, 1743, 1733, 1722,
1711, 1701, 1689, 1679, 1669, 1658, 1648, 1637, 1626, 1616, 1606, 1595, 1585, 1575, 1564, 1554,
1544, 1534, 1524, 1514, 1504, 1494, 1484, 1474, 1464, 1454, 1445, 1435, 1425, 1416, 1406, 1397,
1387, 1378, 1369, 1359, 1350, 1341, 1332, 1323, 1314, 1305, 1296, 1287, 1279, 1270, 1261, 1253),
(2413, 2413, 2412, 2412, 2411, 2410, 2409, 2407, 2406, 2404, 2402, 2399, 2397, 2394, 2391, 2388,
2385, 2381, 2377, 2373, 2369, 2365, 2360, 2355, 2350, 2345, 2340, 2334, 2329, 2323, 2317, 2311,
2304, 2298, 2291, 2284, 2277, 2270, 2263, 2255, 2247, 2240, 2232, 2224, 2216, 2207, 2199, 2190,
2182, 2173, 2164, 2155, 2146, 2137, 2128, 2118, 2109, 2099, 2090, 2080, 2070, 2060, 2051, 2041,
2031, 2020, 2010, 2000, 1990, 1980, 1969, 1959, 1949, 1938, 1927, 1917, 1907, 1896, 1885, 1875,
1865, 1854, 1842, 1833, 1822, 1811, 1801, 1790, 1780, 1769, 1757, 1748, 1737, 1727, 1716, 1705,
1695, 1685, 1674, 1663, 1653, 1643, 1633, 1621, 1612, 1602, 1591, 1581, 1570, 1561, 1551, 1541,
1531, 1521, 1511, 1501, 1491, 1481, 1472, 1462, 1452, 1443, 1433, 1423, 1414, 1405, 1395, 1386,
1377, 1367, 1358, 1349, 1340, 1331, 1322, 1313, 1304, 1296, 1287, 1278, 1270, 1261, 1253, 1244),
(2380, 2380, 2380, 2379, 2379, 2378, 2377, 2375, 2374, 2372, 2370, 2367, 2365, 2362, 2359, 2356,
2353, 2350, 2346, 2342, 2338, 2334, 2329, 2325, 2320, 2315, 2310, 2304, 2299, 2293, 2287, 2281,
2275, 2268, 2262, 2255, 2248, 2241, 2234, 2227, 2219, 2212, 2204, 2196, 2188, 2180, 2172, 2164,
2155, 2147, 2138, 2129, 2121, 2112, 2103, 2093, 2084, 2075, 2066, 2056, 2046, 2037, 2027, 2018,
2008, 1998, 1987, 1978, 1968, 1958, 1948, 1938, 1927, 1917, 1907, 1897, 1887, 1876, 1866, 1856,
1845, 1835, 1824, 1814, 1804, 1793, 1782, 1772, 1762, 1752, 1740, 1731, 1720, 1710, 1700, 1688,
1679, 1669, 1659, 1648, 1637, 1628, 1618, 1608, 1597, 1586, 1577, 1567, 1557, 1547, 1537, 1527,
1518, 1508, 1498, 1488, 1479, 1469, 1459, 1450, 1440, 1431, 1422, 1412, 1403, 1394, 1384, 1375,
1366, 1357, 1348, 1339, 1330, 1321, 1312, 1304, 1295, 1286, 1278, 1269, 1261, 1252, 1244, 1235),
(2349, 2349, 2348, 2348, 2347, 2346, 2345, 2344, 2342, 2340, 2338, 2336, 2334, 2331, 2328, 2325,
2322, 2319, 2315, 2311, 2307, 2303, 2299, 2294, 2290, 2285, 2280, 2275, 2269, 2264, 2258, 2252,
2246, 2240, 2233, 2227, 2220, 2213, 2206, 2199, 2192, 2185, 2177, 2169, 2162, 2154, 2146, 2138,
2129, 2121, 2113, 2104, 2095, 2087, 2078, 2069, 2060, 2051, 2042, 2032, 2023, 2014, 2003, 1995,
1985, 1976, 1966, 1956, 1946, 1935, 1927, 1917, 1907, 1897, 1887, 1876, 1867, 1857, 1846, 1836,
1825, 1816, 1806, 1796, 1785, 1774, 1765, 1755, 1745, 1734, 1723, 1714, 1704, 1694, 1684, 1672,
1663, 1653, 1643, 1633, 1623, 1612, 1603, 1593, 1583, 1573, 1563, 1553, 1544, 1534, 1524, 1514,
1505, 1495, 1485, 1476, 1466, 1457, 1447, 1438, 1429, 1419, 1410, 1401, 1392, 1383, 1374, 1365,
1356, 1347, 1338, 1329, 1320, 1311, 1303, 1294, 1286, 1277, 1269, 1260, 1252, 1243, 1235, 1227),
(2318, 2318, 2317, 2317, 2316, 2315, 2314, 2313, 2311, 2310, 2308, 2305, 2303, 2301, 2298, 2295,
2292, 2289, 2285, 2281, 2278, 2274, 2269, 2265, 2260, 2256, 2251, 2246, 2240, 2235, 2229, 2223,
2218, 2211, 2205, 2199, 2192, 2186, 2179, 2172, 2165, 2158, 2150, 2143, 2135, 2128, 2120, 2112,
2104, 2096, 2087, 2079, 2071, 2062, 2054, 2045, 2036, 2027, 2018, 2009, 2000, 1991, 1982, 1972,
1963, 1953, 1944, 1935, 1925, 1915, 1906, 1896, 1885, 1876, 1867, 1857, 1847, 1837, 1827, 1816,
1807, 1797, 1787, 1777, 1767, 1756, 1747, 1737, 1727, 1717, 1706, 1697, 1687, 1678, 1668, 1658,
1648, 1637, 1628, 1618, 1608, 1598, 1587, 1578, 1569, 1559, 1549, 1540, 1530, 1521, 1511, 1501,
1492, 1482, 1473, 1464, 1454, 1445, 1436, 1426, 1417, 1408, 1399, 1390, 1381, 1372, 1363, 1354,
1345, 1336, 1328, 1319, 1310, 1302, 1293, 1285, 1276, 1268, 1259, 1251, 1243, 1235, 1226, 1218),
(2287, 2287, 2287, 2286, 2286, 2285, 2284, 2282, 2281, 2279, 2277, 2275, 2273, 2271, 2268, 2265,
2262, 2259, 2256, 2252, 2248, 2244, 2240, 2236, 2231, 2227, 2222, 2217, 2212, 2207, 2201, 2195,
2190, 2184, 2178, 2172, 2165, 2159, 2152, 2145, 2138, 2131, 2124, 2117, 2110, 2102, 2094, 2087,
2079, 2071, 2063, 2055, 2046, 2037, 2029, 2020, 2012, 2003, 1995, 1986, 1977, 1968, 1959, 1950,
1941, 1932, 1923, 1913, 1904, 1895, 1884, 1876, 1866, 1857, 1847, 1837, 1828, 1818, 1807, 1799,
1789, 1779, 1769, 1760, 1750, 1739, 1730, 1720, 1711, 1701, 1691, 1680, 1671, 1662, 1652, 1642,
1632, 1623, 1612, 1603, 1593, 1584, 1574, 1565, 1555, 1545, 1536, 1526, 1517, 1507, 1498, 1489,
1479, 1470, 1461, 1451, 1442, 1433, 1424, 1415, 1406, 1397, 1388, 1379, 1370, 1361, 1352, 1344,
1335, 1326, 1318, 1309, 1301, 1292, 1284, 1275, 1267, 1259, 1250, 1242, 1234, 1226, 1218, 1210),
(2258, 2257, 2257, 2257, 2256, 2255, 2254, 2253, 2251, 2250, 2248, 2246, 2244, 2241, 2239, 2236,
2233, 2230, 2227, 2223, 2219, 2216, 2212, 2207, 2203, 2198, 2194, 2189, 2184, 2179, 2173, 2168,
2162, 2157, 2151, 2145, 2138, 2132, 2126, 2119, 2112, 2105, 2098, 2091, 2084, 2077, 2069, 2062,
2054, 2046, 2038, 2031, 2023, 2014, 2006, 1998, 1989, 1981, 1972, 1964, 1955, 1946, 1936, 1929,
1919, 1910, 1901, 1892, 1883, 1874, 1865, 1856, 1846, 1837, 1827, 1818, 1808, 1799, 1790, 1780,
1771, 1761, 1751, 1742, 1731, 1722, 1713, 1703, 1694, 1684, 1675, 1665, 1654, 1646, 1636, 1627,
1617, 1607, 1598, 1587, 1578, 1569, 1560, 1551, 1541, 1532, 1522, 1513, 1504, 1494, 1485, 1476,
1467, 1458, 1448, 1439, 1430, 1421, 1412, 1403, 1394, 1386, 1377, 1368, 1359, 1351, 1342, 1333,
1325, 1316, 1308, 1299, 1291, 1282, 1274, 1266, 1258, 1250, 1241, 1233, 1225, 1217, 1209, 1202),
(2228, 2228, 2228, 2227, 2227, 2226, 2225, 2224, 2222, 2221, 2219, 2217, 2215, 2212, 2210, 2207,
2204, 2201, 2198, 2195, 2191, 2187, 2183, 2179, 2175, 2171, 2166, 2161, 2157, 2152, 2146, 2141,
2136, 2130, 2124, 2118, 2112, 2106, 2100, 2093, 2087, 2080, 2073, 2066, 2059, 2052, 2045, 2037,
2029, 2021, 2015, 2007, 1999, 1991, 1983, 1975, 1967, 1958, 1950, 1942, 1933, 1925, 1916, 1907,
1898, 1890, 1881, 1872, 1863, 1854, 1845, 1836, 1827, 1816, 1807, 1799, 1790, 1780, 1771, 1762,
1753, 1743, 1734, 1723, 1714, 1705, 1696, 1687, 1677, 1668, 1658, 1649, 1640, 1629, 1620, 1611,
1602, 1593, 1583, 1574, 1565, 1555, 1546, 1537, 1527, 1518, 1509, 1500, 1491, 1482, 1472, 1463,
1454, 1445, 1436, 1427, 1419, 1410, 1401, 1392, 1383, 1375, 1366, 1357, 1349, 1340, 1332, 1323,
1315, 1306, 1298, 1290, 1281, 1273, 1265, 1257, 1249, 1241, 1233, 1225, 1217, 1209, 1201, 1193),
(2200, 2200, 2199, 2199, 2198, 2197, 2196, 2195, 2194, 2192, 2190, 2189, 2186, 2184, 2182, 2179,
2176, 2173, 2170, 2167, 2163, 2160, 2156, 2152, 2148, 2144, 2139, 2135, 2130, 2125, 2120, 2115,
2109, 2104, 2098, 2092, 2086, 2080, 2074, 2068, 2062, 2055, 2048, 2042, 2035, 2028, 2020, 2012,
2006, 1999, 1991, 1984, 1976, 1968, 1960, 1952, 1944, 1935, 1927, 1919, 1910, 1902, 1895, 1885,
1878, 1868, 1859, 1851, 1842, 1833, 1824, 1816, 1807, 1798, 1789, 1780, 1771, 1762, 1753, 1744,
1735, 1726, 1716, 1706, 1697, 1688, 1679, 1670, 1661, 1652, 1643, 1633, 1624, 1615, 1606, 1595,
1586, 1578, 1569, 1560, 1550, 1541, 1532, 1523, 1514, 1505, 1496, 1487, 1478, 1469, 1460, 1451,
1442, 1433, 1424, 1416, 1407, 1398, 1389, 1381, 1372, 1364, 1355, 1347, 1338, 1330, 1321, 1313,
1305, 1296, 1288, 1280, 1272, 1264, 1256, 1248, 1240, 1232, 1224, 1216, 1208, 1200, 1193, 1185),
(2172, 2171, 2171, 2171, 2170, 2169, 2168, 2167, 2166, 2164, 2163, 2161, 2159, 2156, 2154, 2152,
2149, 2146, 2143, 2140, 2136, 2133, 2129, 2125, 2121, 2117, 2113, 2108, 2103, 2099, 2094, 2089,
2083, 2078, 2073, 2067, 2061, 2055, 2049, 2043, 2037, 2029, 2024, 2017, 2011, 2003, 1997, 1990,
1983, 1975, 1968, 1961, 1952, 1946, 1938, 1930, 1922, 1914, 1906, 1898, 1890, 1882, 1874, 1865,
1857, 1849, 1840, 1832, 1823, 1814, 1806, 1797, 1788, 1780, 1771, 1762, 1753, 1744, 1735, 1726,
1717, 1708, 1699, 1689, 1680, 1671, 1663, 1654, 1645, 1636, 1627, 1618, 1609, 1600, 1591, 1581,
1572, 1563, 1554, 1545, 1536, 1527, 1518, 1509, 1501, 1492, 1483, 1474, 1465, 1456, 1447, 1439,
1430, 1421, 1413, 1404, 1395, 1387, 1378, 1370, 1361, 1353, 1344, 1336, 1328, 1319, 1311, 1303,
1295, 1286, 1278, 1270, 1262, 1254, 1246, 1238, 1231, 1223, 1215, 1207, 1200, 1192, 1184, 1177),
(2144, 2144, 2144, 2143, 2143, 2142, 2141, 2140, 2138, 2137, 2135, 2133, 2131, 2129, 2127, 2124,
2122, 2119, 2116, 2113, 2110, 2106, 2102, 2099, 2095, 2091, 2086, 2082, 2078, 2073, 2068, 2063,
2058, 2053, 2046, 2042, 2036, 2031, 2025, 2019, 2012, 2006, 2000, 1994, 1986, 1980, 1974, 1967,
1960, 1952, 1944, 1938, 1931, 1923, 1916, 1908, 1901, 1893, 1884, 1876, 1868, 1861, 1853, 1845,
1837, 1829, 1820, 1812, 1804, 1795, 1787, 1778, 1770, 1761, 1752, 1744, 1735, 1726, 1717, 1709,
1700, 1691, 1682, 1672, 1665, 1655, 1646, 1637, 1629, 1620, 1611, 1602, 1593, 1585, 1576, 1567,
1558, 1549, 1540, 1531, 1523, 1514, 1505, 1496, 1487, 1479, 1470, 1461, 1452, 1444, 1435, 1427,
1418, 1409, 1401, 1392, 1384, 1375, 1367, 1359, 1350, 1342, 1334, 1325, 1317, 1309, 1301, 1293,
1285, 1277, 1269, 1261, 1253, 1245, 1237, 1229, 1222, 1214, 1206, 1199, 1191, 1184, 1176, 1169),
(2117, 2117, 2117, 2116, 2116, 2115, 2114, 2113, 2111, 2110, 2108, 2107, 2105, 2103, 2100, 2098,
2095, 2093, 2090, 2087, 2083, 2080, 2076, 2073, 2069, 2065, 2061, 2057, 2052, 2048, 2043, 2037,
2033, 2028, 2023, 2017, 2012, 2006, 2001, 1995, 1989, 1983, 1976, 1969, 1964, 1957, 1951, 1944,
1936, 1930, 1923, 1916, 1909, 1901, 1893, 1887, 1879, 1872, 1864, 1856, 1849, 1841, 1833, 1824,
1816, 1808, 1801, 1793, 1784, 1776, 1768, 1759, 1751, 1743, 1734, 1726, 1717, 1709, 1700, 1691,
1683, 1674, 1666, 1657, 1648, 1640, 1631, 1621, 1612, 1604, 1595, 1586, 1578, 1569, 1561, 1552,
1544, 1535, 1526, 1518, 1509, 1500, 1492, 1483, 1474, 1466, 1457, 1449, 1440, 1431, 1423, 1415,
1406, 1398, 1389, 1381, 1373, 1364, 1356, 1348, 1340, 1331, 1323, 1315, 1307, 1299, 1291, 1283,
1275, 1267, 1259, 1251, 1244, 1236, 1228, 1220, 1213, 1205, 1198, 1190, 1183, 1175, 1168, 1160),
(2090, 2090, 2090, 2090, 2089, 2088, 2087, 2086, 2085, 2084, 2082, 2080, 2078, 2076, 2074, 2072,
2069, 2067, 2064, 2061, 2058, 2054, 2051, 2046, 2044, 2040, 2036, 2031, 2027, 2023, 2018, 2012,
2009, 2003, 1998, 1993, 1987, 1982, 1977, 1970, 1965, 1959, 1952, 1947, 1941, 1934, 1927, 1921,
1915, 1908, 1901, 1893, 1887, 1880, 1873, 1866, 1858, 1850, 1844, 1836, 1828, 1821, 1813, 1805,
1797, 1789, 1782, 1773, 1765, 1756, 1748, 1740, 1733, 1725, 1716, 1708, 1700, 1691, 1683, 1674,
1666, 1658, 1649, 1641, 1632, 1624, 1615, 1606, 1598, 1589, 1581, 1572, 1564, 1555, 1547, 1538,
1529, 1521, 1512, 1504, 1495, 1487, 1478, 1470, 1461, 1453, 1444, 1436, 1428, 1419, 1411, 1403,
1394, 1386, 1378, 1370, 1361, 1353, 1345, 1337, 1329, 1321, 1313, 1305, 1297, 1289, 1281, 1273,
1265, 1258, 1250, 1242, 1234, 1227, 1219, 1212, 1204, 1197, 1189, 1182, 1174, 1167, 1160, 1152),
(2064, 2064, 2064, 2064, 2063, 2062, 2061, 2060, 2059, 2058, 2056, 2055, 2053, 2051, 2049, 2046,
2044, 2041, 2037, 2035, 2032, 2029, 2026, 2021, 2019, 2015, 2011, 2007, 2003, 1998, 1994, 1989,
1984, 1980, 1975, 1969, 1964, 1959, 1952, 1948, 1942, 1935, 1931, 1924, 1918, 1912, 1906, 1899,
1893, 1885, 1880, 1873, 1866, 1859, 1851, 1845, 1838, 1831, 1823, 1816, 1807, 1801, 1793, 1786,
1778, 1770, 1763, 1755, 1747, 1739, 1731, 1722, 1714, 1706, 1699, 1691, 1682, 1674, 1666, 1658,
1649, 1641, 1633, 1625, 1616, 1608, 1599, 1591, 1583, 1574, 1566, 1557, 1549, 1541, 1532, 1524,
1515, 1507, 1499, 1490, 1482, 1474, 1465, 1457, 1449, 1440, 1432, 1424, 1415, 1407, 1399, 1391,
1383, 1375, 1366, 1358, 1350, 1342, 1334, 1326, 1318, 1310, 1302, 1295, 1287, 1279, 1271, 1263,
1256, 1248, 1240, 1233, 1225, 1218, 1210, 1203, 1195, 1188, 1181, 1173, 1166, 1159, 1152, 1145),
(2038, 2038, 2037, 2037, 2037, 2037, 2036, 2035, 2034, 2032, 2031, 2029, 2027, 2025, 2023, 2020,
2019, 2016, 2012, 2011, 2008, 2003, 2001, 1998, 1994, 1990, 1986, 1983, 1978, 1974, 1969, 1965,
1961, 1956, 1951, 1946, 1941, 1935, 1931, 1925, 1919, 1914, 1908, 1901, 1896, 1890, 1884, 1878,
1871, 1865, 1858, 1851, 1845, 1838, 1831, 1824, 1818, 1810, 1803, 1796, 1789, 1781, 1773, 1767,
1759, 1752, 1744, 1736, 1729, 1721, 1713, 1705, 1697, 1688, 1680, 1672, 1665, 1657, 1649, 1641,
1633, 1625, 1617, 1609, 1600, 1592, 1584, 1576, 1568, 1559, 1551, 1543, 1535, 1526, 1518, 1510,
1502, 1493, 1485, 1477, 1469, 1460, 1452, 1444, 1436, 1428, 1420, 1412, 1403, 1395, 1387, 1379,
1371, 1363, 1355, 1347, 1339, 1331, 1323, 1316, 1308, 1300, 1292, 1284, 1277, 1269, 1261, 1254,
1246, 1239, 1231, 1224, 1216, 1209, 1201, 1194, 1187, 1179, 1172, 1165, 1158, 1151, 1144, 1137),
(2014, 2014, 2012, 2012, 2012, 2012, 2011, 2010, 2009, 2007, 2006, 2003, 2003, 2001, 1999, 1995,
1994, 1992, 1989, 1986, 1983, 1980, 1977, 1974, 1969, 1967, 1963, 1959, 1955, 1951, 1947, 1942,
1938, 1933, 1927, 1923, 1918, 1913, 1908, 1902, 1897, 1892, 1885, 1880, 1875, 1868, 1863, 1856,
1850, 1844, 1838, 1831, 1824, 1818, 1811, 1804, 1798, 1790, 1784, 1777, 1769, 1762, 1755, 1748,
1739, 1733, 1726, 1718, 1710, 1703, 1695, 1688, 1680, 1671, 1663, 1655, 1649, 1641, 1633, 1625,
1617, 1609, 1601, 1593, 1585, 1577, 1569, 1561, 1553, 1545, 1537, 1528, 1520, 1512, 1504, 1496,
1488, 1480, 1472, 1464, 1456, 1448, 1440, 1431, 1423, 1415, 1407, 1399, 1391, 1384, 1376, 1368,
1360, 1352, 1344, 1336, 1328, 1321, 1313, 1305, 1297, 1290, 1282, 1274, 1267, 1259, 1252, 1244,
1237, 1229, 1222, 1215, 1207, 1200, 1193, 1185, 1178, 1171, 1164, 1157, 1150, 1143, 1136, 1129),
(1989, 1989, 1989, 1987, 1987, 1986, 1986, 1985, 1984, 1983, 1982, 1980, 1978, 1976, 1974, 1972,
1969, 1968, 1965, 1961, 1959, 1956, 1952, 1950, 1947, 1943, 1939, 1935, 1932, 1927, 1923, 1918,
1915, 1910, 1906, 1901, 1896, 1891, 1885, 1881, 1875, 1870, 1865, 1859, 1853, 1847, 1841, 1836,
1829, 1823, 1816, 1811, 1804, 1798, 1790, 1785, 1778, 1771, 1764, 1756, 1750, 1743, 1736, 1729,
1722, 1714, 1706, 1700, 1693, 1685, 1678, 1670, 1663, 1654, 1646, 1640, 1632, 1624, 1617, 1609,
1601, 1593, 1585, 1578, 1569, 1562, 1554, 1546, 1538, 1530, 1522, 1514, 1506, 1498, 1490, 1482,
1474, 1467, 1459, 1451, 1443, 1435, 1427, 1419, 1411, 1403, 1395, 1387, 1380, 1372, 1364, 1356,
1348, 1341, 1333, 1325, 1318, 1310, 1302, 1295, 1287, 1280, 1272, 1265, 1257, 1250, 1242, 1235,
1227, 1220, 1213, 1206, 1198, 1191, 1184, 1177, 1170, 1163, 1156, 1149, 1142, 1135, 1128, 1121),
(1965, 1965, 1965, 1964, 1964, 1963, 1961, 1961, 1960, 1959, 1958, 1956, 1953, 1952, 1951, 1948,
1946, 1944, 1941, 1939, 1935, 1933, 1930, 1927, 1923, 1919, 1916, 1913, 1909, 1905, 1901, 1897,
1892, 1888, 1883, 1879, 1874, 1868, 1864, 1859, 1854, 1849, 1842, 1838, 1832, 1827, 1821, 1815,
1808, 1803, 1797, 1790, 1784, 1778, 1772, 1765, 1759, 1752, 1745, 1738, 1731, 1725, 1718, 1711,
1704, 1697, 1689, 1682, 1675, 1668, 1660, 1653, 1646, 1637, 1631, 1623, 1616, 1608, 1601, 1593,
1585, 1578, 1569, 1562, 1555, 1547, 1539, 1531, 1524, 1516, 1508, 1500, 1492, 1485, 1477, 1469,
1461, 1453, 1446, 1438, 1430, 1422, 1414, 1407, 1399, 1391, 1383, 1376, 1368, 1360, 1353, 1345,
1337, 1330, 1322, 1315, 1307, 1299, 1292, 1284, 1277, 1270, 1262, 1255, 1247, 1240, 1233, 1225,
1218, 1211, 1204, 1197, 1190, 1182, 1175, 1168, 1161, 1154, 1147, 1141, 1134, 1127, 1120, 1113),
(1941, 1941, 1941, 1940, 1940, 1939, 1939, 1938, 1936, 1935, 1934, 1932, 1931, 1929, 1927, 1925,
1923, 1921, 1918, 1916, 1913, 1910, 1907, 1904, 1901, 1897, 1893, 1890, 1885, 1883, 1879, 1875,
1870, 1866, 1862, 1857, 1851, 1848, 1842, 1838, 1833, 1828, 1822, 1816, 1812, 1806, 1799, 1795,
1789, 1782, 1777, 1771, 1765, 1759, 1752, 1746, 1739, 1733, 1726, 1720, 1713, 1705, 1700, 1693,
1686, 1679, 1671, 1665, 1658, 1651, 1644, 1636, 1629, 1621, 1614, 1607, 1600, 1592, 1585, 1577,
1569, 1562, 1555, 1547, 1540, 1532, 1524, 1517, 1509, 1502, 1494, 1486, 1479, 1471, 1463, 1456,
1448, 1440, 1433, 1425, 1417, 1410, 1402, 1394, 1387, 1379, 1372, 1364, 1356, 1349, 1341, 1334,
1326, 1319, 1311, 1304, 1296, 1289, 1282, 1274, 1267, 1260, 1252, 1245, 1238, 1231, 1223, 1216,
1209, 1202, 1195, 1188, 1181, 1174, 1167, 1160, 1153, 1146, 1139, 1132, 1126, 1119, 1112, 1106),
(1918, 1918, 1918, 1917, 1917, 1916, 1915, 1914, 1913, 1912, 1910, 1909, 1908, 1906, 1904, 1901,
1900, 1898, 1895, 1893, 1890, 1887, 1884, 1881, 1878, 1875, 1872, 1867, 1864, 1861, 1857, 1853,
1849, 1844, 1840, 1836, 1831, 1827, 1822, 1816, 1812, 1807, 1802, 1797, 1790, 1786, 1780, 1774,
1769, 1763, 1756, 1751, 1745, 1739, 1733, 1727, 1721, 1714, 1708, 1702, 1695, 1688, 1682, 1675,
1668, 1661, 1654, 1648, 1641, 1634, 1627, 1620, 1612, 1604, 1598, 1591, 1584, 1577, 1569, 1562,
1555, 1547, 1540, 1532, 1525, 1517, 1510, 1503, 1495, 1488, 1480, 1473, 1465, 1458, 1450, 1442,
1435, 1427, 1420, 1412, 1405, 1397, 1390, 1382, 1375, 1367, 1360, 1352, 1345, 1338, 1330, 1323,
1315, 1308, 1301, 1293, 1286, 1279, 1271, 1264, 1257, 1250, 1243, 1235, 1228, 1221, 1214, 1207,
1200, 1193, 1186, 1179, 1172, 1165, 1158, 1152, 1145, 1138, 1131, 1125, 1118, 1111, 1105, 1098),
(1895, 1895, 1895, 1893, 1893, 1893, 1892, 1892, 1891, 1889, 1888, 1887, 1884, 1883, 1882, 1880,
1878, 1875, 1873, 1871, 1867, 1865, 1862, 1859, 1856, 1853, 1850, 1846, 1842, 1839, 1835, 1831,
1827, 1823, 1819, 1815, 1810, 1806, 1801, 1796, 1791, 1787, 1782, 1776, 1771, 1765, 1761, 1755,
1748, 1744, 1738, 1731, 1726, 1721, 1714, 1708, 1702, 1696, 1689, 1683, 1677, 1671, 1663, 1658,
1651, 1644, 1637, 1631, 1624, 1617, 1610, 1603, 1595, 1589, 1582, 1575, 1568, 1561, 1554, 1547,
1539, 1532, 1525, 1518, 1510, 1503, 1496, 1488, 1481, 1474, 1466, 1459, 1452, 1444, 1437, 1429,
1422, 1415, 1407, 1400, 1393, 1385, 1378, 1370, 1363, 1356, 1348, 1341, 1334, 1326, 1319, 1312,
1305, 1297, 1290, 1283, 1276, 1268, 1261, 1254, 1247, 1240, 1233, 1226, 1219, 1212, 1205, 1198,
1191, 1184, 1177, 1170, 1164, 1157, 1150, 1143, 1137, 1130, 1123, 1117, 1110, 1103, 1097, 1090),
(1872, 1872, 1872, 1872, 1871, 1871, 1870, 1868, 1867, 1867, 1866, 1864, 1863, 1861, 1859, 1858,
1855, 1853, 1850, 1849, 1846, 1842, 1841, 1838, 1835, 1832, 1828, 1824, 1822, 1818, 1814, 1810,
1806, 1802, 1798, 1794, 1790, 1785, 1781, 1776, 1771, 1767, 1762, 1756, 1752, 1746, 1740, 1736,
1730, 1725, 1719, 1714, 1708, 1702, 1696, 1689, 1684, 1678, 1671, 1666, 1659, 1653, 1646, 1640,
1634, 1627, 1620, 1614, 1607, 1601, 1594, 1586, 1580, 1574, 1567, 1560, 1553, 1546, 1539, 1532,
1525, 1517, 1510, 1503, 1496, 1489, 1482, 1475, 1467, 1460, 1453, 1446, 1438, 1431, 1424, 1417,
1409, 1402, 1395, 1388, 1380, 1373, 1366, 1359, 1351, 1344, 1337, 1330, 1323, 1315, 1308, 1301,
1294, 1287, 1280, 1273, 1265, 1258, 1251, 1244, 1237, 1230, 1223, 1216, 1209, 1203, 1196, 1189,
1182, 1175, 1168, 1162, 1155, 1148, 1142, 1135, 1128, 1122, 1115, 1109, 1102, 1096, 1089, 1083),
(1850, 1850, 1850, 1850, 1849, 1849, 1848, 1847, 1846, 1845, 1844, 1842, 1841, 1839, 1838, 1836,
1833, 1832, 1829, 1827, 1824, 1822, 1819, 1816, 1814, 1810, 1807, 1804, 1801, 1797, 1793, 1790,
1786, 1782, 1778, 1773, 1770, 1765, 1761, 1756, 1752, 1747, 1742, 1737, 1731, 1727, 1722, 1717,
1711, 1705, 1701, 1695, 1688, 1684, 1678, 1671, 1666, 1660, 1654, 1648, 1642, 1636, 1629, 1623,
1617, 1611, 1603, 1598, 1591, 1585, 1578, 1570, 1565, 1558, 1551, 1544, 1537, 1531, 1524, 1517,
1510, 1503, 1496, 1489, 1482, 1475, 1468, 1461, 1454, 1447, 1440, 1432, 1425, 1418, 1411, 1404,
1397, 1390, 1383, 1375, 1368, 1361, 1354, 1347, 1340, 1333, 1326, 1319, 1311, 1304, 1297, 1290,
1283, 1276, 1269, 1262, 1255, 1248, 1241, 1234, 1228, 1221, 1214, 1207, 1200, 1193, 1187, 1180,
1173, 1166, 1160, 1153, 1147, 1140, 1133, 1127, 1120, 1114, 1107, 1101, 1095, 1088, 1082, 1076),
(1829, 1829, 1828, 1828, 1828, 1827, 1825, 1825, 1824, 1823, 1822, 1821, 1819, 1818, 1816, 1814,
1812, 1810, 1807, 1806, 1804, 1801, 1798, 1796, 1793, 1790, 1787, 1782, 1780, 1777, 1773, 1769,
1765, 1762, 1757, 1754, 1750, 1745, 1740, 1737, 1731, 1728, 1722, 1718, 1713, 1708, 1703, 1697,
1693, 1688, 1682, 1677, 1671, 1666, 1660, 1654, 1649, 1643, 1637, 1631, 1625, 1619, 1612, 1607,
1600, 1594, 1587, 1581, 1575, 1569, 1562, 1556, 1549, 1542, 1536, 1529, 1522, 1516, 1509, 1502,
1495, 1489, 1482, 1475, 1468, 1461, 1454, 1447, 1440, 1433, 1426, 1419, 1412, 1405, 1398, 1391,
1384, 1377, 1370, 1363, 1356, 1349, 1342, 1335, 1328, 1321, 1314, 1307, 1301, 1294, 1287, 1280,
1273, 1266, 1259, 1252, 1245, 1238, 1232, 1225, 1218, 1211, 1204, 1198, 1191, 1184, 1178, 1171,
1164, 1158, 1151, 1145, 1138, 1132, 1125, 1119, 1112, 1106, 1100, 1093, 1087, 1081, 1074, 1068),
(1807, 1807, 1807, 1807, 1806, 1806, 1805, 1804, 1803, 1802, 1801, 1799, 1798, 1797, 1795, 1793,
1791, 1790, 1787, 1785, 1782, 1780, 1778, 1774, 1772, 1769, 1765, 1763, 1760, 1756, 1753, 1748,
1746, 1742, 1738, 1734, 1730, 1726, 1722, 1717, 1713, 1708, 1704, 1699, 1694, 1689, 1685, 1680,
1675, 1669, 1663, 1659, 1653, 1648, 1642, 1637, 1631, 1626, 1620, 1614, 1608, 1602, 1595, 1590,
1584, 1578, 1572, 1565, 1559, 1553, 1547, 1540, 1534, 1527, 1521, 1514, 1508, 1501, 1494, 1488,
1481, 1474, 1468, 1461, 1454, 1447, 1441, 1434, 1427, 1420, 1413, 1407, 1400, 1393, 1386, 1379,
1372, 1365, 1358, 1352, 1345, 1338, 1331, 1324, 1317, 1310, 1303, 1297, 1290, 1283, 1276, 1269,
1262, 1256, 1249, 1242, 1235, 1229, 1222, 1215, 1209, 1202, 1195, 1189, 1182, 1175, 1169, 1162,
1156, 1149, 1143, 1136, 1130, 1123, 1117, 1111, 1104, 1098, 1092, 1086, 1079, 1073, 1067, 1061),
(1786, 1786, 1786, 1786, 1785, 1785, 1784, 1782, 1782, 1781, 1780, 1779, 1778, 1776, 1774, 1773,
1771, 1769, 1767, 1765, 1762, 1760, 1756, 1755, 1752, 1748, 1746, 1743, 1739, 1737, 1733, 1730,
1726, 1722, 1719, 1714, 1711, 1706, 1703, 1697, 1694, 1689, 1685, 1680, 1676, 1671, 1666, 1662,
1657, 1651, 1646, 1641, 1636, 1631, 1625, 1620, 1614, 1609, 1603, 1597, 1591, 1586, 1580, 1574,
1568, 1562, 1556, 1550, 1544, 1537, 1531, 1525, 1519, 1512, 1506, 1499, 1493, 1487, 1480, 1474,
1467, 1460, 1454, 1447, 1441, 1434, 1427, 1421, 1414, 1407, 1401, 1394, 1387, 1380, 1374, 1367,
1360, 1353, 1347, 1340, 1333, 1326, 1319, 1313, 1306, 1299, 1292, 1286, 1279, 1272, 1266, 1259,
1252, 1245, 1239, 1232, 1226, 1219, 1212, 1206, 1199, 1193, 1186, 1179, 1173, 1166, 1160, 1154,
1147, 1141, 1134, 1128, 1122, 1115, 1109, 1103, 1097, 1090, 1084, 1078, 1072, 1066, 1060, 1054),
(1765, 1765, 1765, 1765, 1765, 1764, 1764, 1763, 1762, 1761, 1760, 1759, 1756, 1756, 1754, 1752,
1751, 1748, 1747, 1745, 1742, 1739, 1737, 1735, 1731, 1729, 1727, 1723, 1720, 1717, 1714, 1710,
1706, 1703, 1700, 1696, 1692, 1688, 1684, 1680, 1676, 1671, 1667, 1662, 1658, 1653, 1648, 1644,
1638, 1634, 1629, 1624, 1619, 1612, 1608, 1603, 1597, 1592, 1586, 1581, 1575, 1569, 1564, 1558,
1552, 1546, 1540, 1534, 1528, 1522, 1516, 1510, 1504, 1497, 1491, 1485, 1479, 1472, 1466, 1460,
1453, 1447, 1440, 1434, 1427, 1421, 1414, 1408, 1401, 1394, 1388, 1381, 1375, 1368, 1361, 1355,
1348, 1341, 1335, 1328, 1321, 1315, 1308, 1302, 1295, 1288, 1282, 1275, 1268, 1262, 1255, 1249,
1242, 1235, 1229, 1222, 1216, 1209, 1203, 1196, 1190, 1183, 1177, 1170, 1164, 1158, 1151, 1145,
1139, 1132, 1126, 1120, 1114, 1107, 1101, 1095, 1089, 1083, 1077, 1070, 1064, 1058, 1052, 1046),
(1746, 1745, 1745, 1745, 1745, 1744, 1743, 1743, 1742, 1740, 1739, 1739, 1737, 1736, 1734, 1733,
1731, 1729, 1727, 1725, 1722, 1720, 1718, 1714, 1713, 1710, 1706, 1704, 1701, 1697, 1695, 1691,
1688, 1685, 1680, 1677, 1672, 1670, 1666, 1662, 1657, 1653, 1649, 1644, 1640, 1635, 1631, 1626,
1620, 1617, 1612, 1607, 1602, 1595, 1591, 1586, 1581, 1575, 1569, 1565, 1559, 1553, 1548, 1542,
1536, 1531, 1525, 1519, 1513, 1507, 1501, 1495, 1489, 1483, 1477, 1471, 1464, 1458, 1452, 1446,
1439, 1433, 1427, 1420, 1414, 1408, 1401, 1395, 1388, 1382, 1375, 1369, 1362, 1356, 1349, 1343,
1336, 1330, 1323, 1317, 1310, 1304, 1297, 1291, 1284, 1277, 1271, 1264, 1258, 1251, 1245, 1238,
1232, 1225, 1219, 1213, 1206, 1200, 1193, 1187, 1181, 1174, 1168, 1162, 1155, 1149, 1143, 1136,
1130, 1124, 1118, 1112, 1105, 1099, 1093, 1087, 1081, 1075, 1069, 1063, 1057, 1051, 1045, 1039),
(1726, 1726, 1725, 1725, 1725, 1723, 1723, 1722, 1722, 1721, 1720, 1719, 1717, 1716, 1714, 1713,
1711, 1709, 1706, 1705, 1703, 1701, 1699, 1696, 1694, 1691, 1688, 1685, 1682, 1679, 1676, 1672,
1669, 1666, 1662, 1659, 1654, 1651, 1646, 1643, 1638, 1635, 1631, 1627, 1621, 1618, 1612, 1609,
1603, 1599, 1595, 1590, 1585, 1580, 1575, 1569, 1564, 1559, 1554, 1549, 1543, 1538, 1532, 1527,
1521, 1515, 1510, 1504, 1498, 1492, 1486, 1480, 1474, 1469, 1463, 1456, 1450, 1444, 1438, 1432,
1426, 1420, 1413, 1407, 1401, 1395, 1388, 1382, 1376, 1369, 1363, 1357, 1350, 1344, 1337, 1331,
1325, 1318, 1312, 1305, 1299, 1292, 1286, 1280, 1273, 1267, 1260, 1254, 1248, 1241, 1235, 1228,
1222, 1216, 1209, 1203, 1197, 1190, 1184, 1178, 1171, 1165, 1159, 1153, 1146, 1140, 1134, 1128,
1122, 1116, 1110, 1103, 1097, 1091, 1085, 1079, 1073, 1067, 1061, 1056, 1050, 1044, 1038, 1032),
(1705, 1705, 1705, 1705, 1705, 1705, 1704, 1703, 1703, 1702, 1701, 1699, 1697, 1697, 1695, 1694,
1692, 1689, 1688, 1686, 1684, 1682, 1680, 1677, 1675, 1671, 1669, 1667, 1663, 1661, 1658, 1654,
1651, 1648, 1644, 1641, 1637, 1633, 1629, 1626, 1621, 1618, 1614, 1609, 1604, 1601, 1595, 1592,
1586, 1583, 1578, 1573, 1568, 1563, 1558, 1553, 1548, 1543, 1538, 1533, 1527, 1522, 1517, 1511,
1506, 1500, 1495, 1489, 1483, 1478, 1472, 1466, 1460, 1454, 1448, 1443, 1437, 1431, 1425, 1419,
1412, 1406, 1400, 1394, 1388, 1382, 1376, 1369, 1363, 1357, 1351, 1344, 1338, 1332, 1326, 1319,
1313, 1307, 1300, 1294, 1288, 1281, 1275, 1269, 1263, 1256, 1250, 1244, 1237, 1231, 1225, 1218,
1212, 1206, 1200, 1193, 1187, 1181, 1175, 1169, 1162, 1156, 1150, 1144, 1138, 1132, 1126, 1120,
1113, 1107, 1101, 1095, 1089, 1084, 1078, 1072, 1066, 1060, 1054, 1048, 1042, 1037, 1031, 1025),
(1687, 1687, 1687, 1686, 1686, 1685, 1685, 1684, 1683, 1682, 1680, 1680, 1679, 1678, 1676, 1675,
1672, 1671, 1669, 1668, 1665, 1663, 1661, 1659, 1655, 1654, 1651, 1648, 1645, 1642, 1638, 1636,
1633, 1629, 1626, 1623, 1619, 1616, 1612, 1608, 1603, 1600, 1595, 1592, 1587, 1584, 1580, 1575,
1570, 1566, 1561, 1557, 1552, 1547, 1542, 1537, 1533, 1527, 1522, 1517, 1512, 1507, 1501, 1496,
1491, 1485, 1480, 1474, 1469, 1463, 1457, 1452, 1446, 1440, 1435, 1429, 1423, 1417, 1411, 1405,
1399, 1393, 1387, 1381, 1375, 1369, 1363, 1357, 1351, 1345, 1339, 1332, 1326, 1320, 1314, 1308,
1302, 1295, 1289, 1283, 1277, 1271, 1264, 1258, 1252, 1246, 1240, 1233, 1227, 1221, 1215, 1209,
1202, 1196, 1190, 1184, 1178, 1172, 1166, 1160, 1153, 1147, 1141, 1135, 1129, 1123, 1117, 1111,
1105, 1099, 1093, 1087, 1082, 1076, 1070, 1064, 1058, 1052, 1047, 1041, 1035, 1030, 1024, 1018),
(1668, 1668, 1668, 1667, 1667, 1667, 1666, 1665, 1665, 1663, 1663, 1662, 1660, 1659, 1658, 1655,
1654, 1653, 1651, 1649, 1646, 1645, 1643, 1640, 1637, 1635, 1633, 1629, 1627, 1625, 1621, 1619,
1615, 1612, 1609, 1604, 1602, 1598, 1595, 1591, 1586, 1583, 1578, 1575, 1570, 1567, 1563, 1559,
1554, 1550, 1545, 1541, 1536, 1531, 1527, 1522, 1517, 1512, 1507, 1502, 1497, 1492, 1486, 1481,
1476, 1471, 1465, 1460, 1454, 1449, 1443, 1438, 1432, 1427, 1421, 1415, 1409, 1404, 1398, 1392,
1386, 1380, 1374, 1369, 1363, 1357, 1351, 1345, 1339, 1333, 1327, 1321, 1315, 1309, 1302, 1296,
1290, 1284, 1278, 1272, 1266, 1260, 1254, 1248, 1242, 1235, 1229, 1223, 1217, 1211, 1205, 1199,
1193, 1187, 1181, 1175, 1169, 1163, 1157, 1151, 1145, 1139, 1133, 1127, 1121, 1115, 1109, 1103,
1097, 1091, 1085, 1080, 1074, 1068, 1062, 1057, 1051, 1045, 1039, 1034, 1028, 1022, 1017, 1010),
(1649, 1649, 1649, 1649, 1649, 1648, 1646, 1646, 1646, 1645, 1644, 1643, 1642, 1641, 1638, 1637,
1636, 1635, 1633, 1631, 1629, 1627, 1625, 1621, 1620, 1618, 1615, 1612, 1610, 1607, 1603, 1601,
1598, 1595, 1592, 1587, 1585, 1581, 1578, 1574, 1569, 1567, 1563, 1559, 1555, 1551, 1547, 1542,
1538, 1534, 1529, 1525, 1520, 1516, 1511, 1506, 1501, 1497, 1492, 1487, 1482, 1477, 1472, 1467,
1461, 1456, 1451, 1446, 1440, 1435, 1429, 1424, 1418, 1413, 1407, 1402, 1396, 1390, 1385, 1379,
1373, 1368, 1362, 1356, 1350, 1344, 1338, 1333, 1327, 1321, 1315, 1309, 1303, 1297, 1291, 1285,
1279, 1273, 1267, 1261, 1255, 1249, 1243, 1237, 1231, 1225, 1219, 1213, 1207, 1201, 1195, 1189,
1183, 1177, 1171, 1165, 1159, 1154, 1148, 1142, 1136, 1130, 1124, 1118, 1112, 1106, 1101, 1095,
1089, 1083, 1078, 1072, 1066, 1060, 1055, 1049, 1043, 1038, 1032, 1027, 1021, 1014, 1010, 1004),
(1631, 1631, 1631, 1631, 1629, 1629, 1629, 1629, 1628, 1627, 1626, 1625, 1624, 1623, 1620, 1620,
1618, 1617, 1615, 1612, 1611, 1609, 1607, 1604, 1602, 1600, 1598, 1595, 1592, 1590, 1586, 1584,
1581, 1578, 1575, 1570, 1568, 1565, 1561, 1558, 1554, 1550, 1546, 1543, 1539, 1535, 1531, 1526,
1522, 1518, 1514, 1509, 1505, 1500, 1496, 1491, 1486, 1482, 1477, 1472, 1467, 1462, 1457, 1452,
1447, 1442, 1437, 1432, 1426, 1421, 1416, 1410, 1405, 1399, 1394, 1389, 1383, 1377, 1372, 1366,
1361, 1355, 1349, 1344, 1338, 1332, 1326, 1321, 1315, 1309, 1303, 1297, 1292, 1286, 1280, 1274,
1268, 1262, 1256, 1250, 1245, 1239, 1233, 1227, 1221, 1215, 1209, 1203, 1197, 1191, 1186, 1180,
1174, 1168, 1162, 1156, 1150, 1145, 1139, 1133, 1127, 1121, 1115, 1110, 1104, 1098, 1092, 1087,
1081, 1075, 1070, 1064, 1058, 1053, 1047, 1042, 1036, 1030, 1025, 1018, 1014, 1008, 1003, 997),
(1612, 1612, 1612, 1612, 1612, 1612, 1611, 1611, 1610, 1609, 1608, 1607, 1606, 1604, 1603, 1602,
1601, 1599, 1597, 1595, 1594, 1592, 1589, 1586, 1585, 1583, 1580, 1578, 1575, 1572, 1569, 1567,
1564, 1561, 1558, 1555, 1551, 1548, 1545, 1541, 1538, 1534, 1530, 1526, 1523, 1519, 1515, 1511,
1507, 1502, 1498, 1494, 1489, 1485, 1481, 1476, 1471, 1467, 1462, 1457, 1453, 1448, 1443, 1438,
1433, 1428, 1423, 1418, 1413, 1407, 1402, 1397, 1392, 1386, 1381, 1375, 1370, 1365, 1359, 1354,
1348, 1343, 1337, 1331, 1326, 1320, 1315, 1309, 1303, 1297, 1292, 1286, 1280, 1275, 1269, 1263,
1257, 1251, 1246, 1240, 1234, 1228, 1222, 1217, 1211, 1205, 1199, 1193, 1188, 1182, 1176, 1170,
1164, 1159, 1153, 1147, 1141, 1136, 1130, 1124, 1118, 1113, 1107, 1101, 1096, 1090, 1084, 1079,
1073, 1068, 1062, 1056, 1051, 1045, 1040, 1034, 1029, 1023, 1018, 1012, 1007, 1001, 996, 991),
(1595, 1595, 1595, 1595, 1595, 1594, 1594, 1593, 1592, 1592, 1591, 1590, 1587, 1586, 1586, 1585,
1583, 1582, 1580, 1578, 1576, 1574, 1572, 1569, 1568, 1566, 1563, 1561, 1558, 1556, 1553, 1550,
1547, 1544, 1541, 1538, 1535, 1532, 1528, 1525, 1521, 1518, 1514, 1511, 1507, 1503, 1499, 1495,
1491, 1487, 1483, 1479, 1474, 1470, 1466, 1461, 1457, 1452, 1448, 1443, 1438, 1433, 1429, 1424,
1419, 1414, 1409, 1404, 1399, 1394, 1389, 1384, 1378, 1373, 1368, 1363, 1357, 1352, 1347, 1341,
1336, 1330, 1325, 1319, 1314, 1308, 1303, 1297, 1292, 1286, 1280, 1275, 1269, 1263, 1258, 1252,
1246, 1241, 1235, 1229, 1224, 1218, 1212, 1207, 1201, 1195, 1189, 1184, 1178, 1172, 1167, 1161,
1155, 1150, 1144, 1138, 1133, 1127, 1121, 1116, 1110, 1104, 1099, 1093, 1088, 1082, 1076, 1071,
1065, 1060, 1054, 1049, 1043, 1038, 1032, 1027, 1022, 1016, 1010, 1005, 1000, 995, 989, 984),
(1578, 1578, 1578, 1578, 1577, 1577, 1576, 1576, 1575, 1574, 1573, 1572, 1570, 1569, 1569, 1567,
1566, 1564, 1563, 1561, 1559, 1557, 1555, 1553, 1551, 1549, 1547, 1544, 1542, 1539, 1536, 1534,
1531, 1528, 1525, 1522, 1519, 1516, 1512, 1509, 1506, 1502, 1499, 1495, 1491, 1488, 1484, 1480,
1476, 1472, 1468, 1464, 1459, 1455, 1451, 1447, 1442, 1438, 1433, 1429, 1424, 1419, 1415, 1410,
1405, 1400, 1395, 1391, 1386, 1381, 1376, 1370, 1365, 1360, 1355, 1350, 1345, 1339, 1334, 1329,
1324, 1318, 1313, 1307, 1302, 1297, 1291, 1286, 1280, 1275, 1269, 1264, 1258, 1253, 1247, 1241,
1236, 1230, 1225, 1219, 1213, 1208, 1202, 1197, 1191, 1185, 1180, 1174, 1169, 1163, 1157, 1152,
1146, 1141, 1135, 1129, 1124, 1118, 1113, 1107, 1102, 1096, 1090, 1085, 1079, 1074, 1068, 1063,
1058, 1052, 1047, 1041, 1036, 1030, 1025, 1020, 1014, 1009, 1004, 997, 993, 988, 983, 978),
(1561, 1561, 1561, 1561, 1560, 1560, 1559, 1559, 1558, 1557, 1556, 1555, 1554, 1553, 1552, 1551,
1549, 1548, 1546, 1544, 1543, 1541, 1539, 1537, 1535, 1532, 1530, 1528, 1525, 1523, 1520, 1518,
1515, 1512, 1509, 1506, 1503, 1500, 1497, 1493, 1490, 1487, 1483, 1480, 1476, 1472, 1469, 1465,
1461, 1457, 1453, 1449, 1445, 1441, 1436, 1432, 1428, 1423, 1419, 1415, 1410, 1406, 1401, 1396,
1392, 1387, 1382, 1377, 1372, 1367, 1363, 1358, 1353, 1348, 1342, 1337, 1332, 1327, 1322, 1317,
1311, 1306, 1301, 1296, 1290, 1285, 1280, 1274, 1269, 1264, 1258, 1253, 1247, 1242, 1236, 1231,
1225, 1220, 1214, 1209, 1203, 1198, 1192, 1187, 1181, 1176, 1170, 1165, 1159, 1154, 1148, 1143,
1137, 1132, 1126, 1121, 1115, 1110, 1104, 1099, 1093, 1088, 1082, 1077, 1071, 1066, 1061, 1055,
1050, 1044, 1039, 1034, 1028, 1023, 1018, 1013, 1007, 1001, 997, 992, 986, 980, 976, 971),
(1544, 1544, 1544, 1544, 1543, 1543, 1542, 1542, 1541, 1540, 1540, 1539, 1538, 1536, 1535, 1534,
1533, 1531, 1530, 1528, 1526, 1524, 1522, 1520, 1518, 1516, 1514, 1512, 1509, 1507, 1504, 1502,
1499, 1496, 1493, 1490, 1487, 1484, 1481, 1478, 1475, 1471, 1468, 1465, 1461, 1457, 1454, 1450,
1446, 1442, 1438, 1434, 1430, 1426, 1422, 1418, 1414, 1409, 1405, 1401, 1396, 1392, 1387, 1383,
1378, 1374, 1369, 1364, 1359, 1355, 1350, 1345, 1340, 1335, 1330, 1325, 1320, 1315, 1310, 1305,
1300, 1294, 1289, 1284, 1279, 1274, 1268, 1263, 1258, 1252, 1247, 1242, 1236, 1231, 1226, 1220,
1215, 1210, 1204, 1199, 1193, 1188, 1182, 1177, 1172, 1166, 1161, 1155, 1150, 1144, 1139, 1134,
1128, 1123, 1117, 1112, 1106, 1101, 1096, 1090, 1085, 1079, 1074, 1069, 1063, 1058, 1053, 1047,
1042, 1037, 1032, 1026, 1021, 1016, 1010, 1005, 1000, 995, 990, 984, 980, 975, 969, 963),
(1528, 1528, 1527, 1527, 1527, 1526, 1526, 1525, 1525, 1524, 1523, 1522, 1521, 1520, 1519, 1518,
1516, 1515, 1513, 1512, 1510, 1508, 1506, 1504, 1502, 1500, 1498, 1496, 1493, 1491, 1489, 1486,
1483, 1481, 1478, 1475, 1472, 1469, 1466, 1463, 1460, 1456, 1453, 1450, 1446, 1443, 1439, 1435,
1432, 1428, 1424, 1420, 1416, 1412, 1408, 1404, 1400, 1396, 1391, 1387, 1383, 1378, 1374, 1369,
1365, 1360, 1356, 1351, 1346, 1342, 1337, 1332, 1327, 1323, 1318, 1313, 1308, 1303, 1298, 1293,
1288, 1283, 1278, 1273, 1267, 1262, 1257, 1252, 1247, 1242, 1236, 1231, 1226, 1221, 1215, 1210,
1205, 1199, 1194, 1189, 1183, 1178, 1173, 1167, 1162, 1157, 1151, 1146, 1141, 1135, 1130, 1125,
1119, 1114, 1109, 1103, 1098, 1093, 1087, 1082, 1077, 1071, 1066, 1061, 1056, 1050, 1045, 1040,
1035, 1029, 1024, 1018, 1014, 1009, 1004, 997, 993, 988, 983, 978, 973, 967, 963, 958),
(1511, 1511, 1511, 1511, 1511, 1510, 1510, 1509, 1508, 1508, 1507, 1506, 1505, 1504, 1503, 1502,
1500, 1499, 1497, 1496, 1494, 1492, 1491, 1489, 1487, 1485, 1482, 1480, 1478, 1476, 1473, 1471,
1468, 1465, 1463, 1460, 1457, 1454, 1451, 1448, 1445, 1442, 1438, 1435, 1432, 1428, 1425, 1421,
1417, 1414, 1410, 1406, 1402, 1398, 1394, 1390, 1386, 1382, 1378, 1374, 1369, 1365, 1361, 1356,
1352, 1347, 1343, 1338, 1334, 1329, 1325, 1320, 1315, 1310, 1306, 1301, 1296, 1291, 1286, 1281,
1276, 1271, 1266, 1261, 1256, 1251, 1246, 1241, 1236, 1231, 1226, 1220, 1215, 1210, 1205, 1200,
1195, 1189, 1184, 1179, 1174, 1168, 1163, 1158, 1153, 1147, 1142, 1137, 1132, 1126, 1121, 1116,
1110, 1105, 1100, 1095, 1089, 1084, 1079, 1074, 1069, 1063, 1058, 1053, 1048, 1043, 1037, 1032,
1027, 1022, 1017, 1012, 1007, 1001, 996, 991, 986, 980, 976, 971, 966, 961, 956, 950),
(1495, 1495, 1495, 1495, 1495, 1494, 1494, 1493, 1493, 1492, 1491, 1490, 1489, 1488, 1487, 1486,
1484, 1483, 1482, 1480, 1478, 1477, 1475, 1473, 1471, 1469, 1467, 1465, 1463, 1460, 1458, 1455,
1453, 1450, 1448, 1445, 1442, 1439, 1436, 1433, 1430, 1427, 1424, 1420, 1417, 1414, 1410, 1407,
1403, 1400, 1396, 1392, 1388, 1385, 1381, 1377, 1373, 1369, 1365, 1360, 1356, 1352, 1348, 1343,
1339, 1335, 1330, 1326, 1321, 1317, 1312, 1308, 1303, 1298, 1294, 1289, 1284, 1279, 1274, 1270,
1265, 1260, 1255, 1250, 1245, 1240, 1235, 1230, 1225, 1220, 1215, 1210, 1205, 1200, 1195, 1190,
1184, 1179, 1174, 1169, 1164, 1159, 1154, 1148, 1143, 1138, 1133, 1128, 1123, 1117, 1112, 1107,
1102, 1097, 1091, 1086, 1081, 1076, 1071, 1066, 1060, 1055, 1050, 1045, 1040, 1035, 1030, 1025,
1020, 1014, 1010, 1005, 999, 993, 989, 984, 979, 975, 970, 965, 959, 955, 950, 945),
(1479, 1479, 1479, 1479, 1479, 1478, 1478, 1477, 1477, 1476, 1475, 1474, 1473, 1472, 1471, 1470,
1469, 1467, 1466, 1465, 1463, 1461, 1460, 1458, 1456, 1454, 1452, 1450, 1447, 1445, 1443, 1440,
1438, 1435, 1433, 1430, 1427, 1425, 1422, 1419, 1416, 1413, 1409, 1406, 1403, 1400, 1396, 1393,
1389, 1386, 1382, 1378, 1375, 1371, 1367, 1363, 1359, 1355, 1351, 1347, 1343, 1339, 1335, 1331,
1326, 1322, 1318, 1313, 1309, 1305, 1300, 1295, 1291, 1286, 1282, 1277, 1272, 1268, 1263, 1258,
1253, 1249, 1244, 1239, 1234, 1229, 1224, 1219, 1215, 1210, 1205, 1200, 1195, 1190, 1185, 1180,
1175, 1170, 1164, 1159, 1154, 1149, 1144, 1139, 1134, 1129, 1124, 1119, 1114, 1108, 1103, 1098,
1093, 1088, 1083, 1078, 1073, 1068, 1063, 1058, 1053, 1047, 1042, 1037, 1032, 1027, 1022, 1017,
1012, 1007, 1001, 997, 992, 987, 983, 978, 973, 967, 963, 958, 953, 948, 944, 939),
(1464, 1464, 1464, 1464, 1463, 1463, 1462, 1462, 1461, 1461, 1460, 1459, 1458, 1457, 1456, 1455,
1454, 1452, 1451, 1449, 1448, 1446, 1444, 1443, 1441, 1439, 1437, 1435, 1433, 1430, 1428, 1426,
1423, 1421, 1418, 1416, 1413, 1410, 1407, 1404, 1401, 1398, 1395, 1392, 1389, 1386, 1382, 1379,
1376, 1372, 1369, 1365, 1361, 1358, 1354, 1350, 1346, 1342, 1338, 1334, 1330, 1326, 1322, 1318,
1314, 1310, 1305, 1301, 1297, 1292, 1288, 1284, 1279, 1275, 1270, 1266, 1261, 1256, 1252, 1247,
1242, 1238, 1233, 1228, 1223, 1219, 1214, 1209, 1204, 1199, 1194, 1189, 1184, 1180, 1175, 1170,
1165, 1160, 1155, 1150, 1145, 1140, 1135, 1130, 1125, 1120, 1115, 1110, 1105, 1100, 1095, 1090,
1085, 1080, 1075, 1070, 1065, 1060, 1055, 1050, 1045, 1040, 1035, 1030, 1025, 1020, 1014, 1010,
1005, 1000, 995, 990, 984, 980, 976, 971, 966, 961, 956, 952, 946, 942, 937, 932),
(1449, 1449, 1448, 1448, 1448, 1448, 1447, 1447, 1446, 1445, 1445, 1444, 1443, 1442, 1441, 1440,
1438, 1437, 1436, 1434, 1433, 1431, 1430, 1428, 1426, 1424, 1422, 1420, 1418, 1416, 1414, 1411,
1409, 1406, 1404, 1401, 1399, 1396, 1393, 1390, 1387, 1384, 1381, 1378, 1375, 1372, 1369, 1365,
1362, 1359, 1355, 1352, 1348, 1344, 1341, 1337, 1333, 1329, 1326, 1322, 1318, 1314, 1310, 1306,
1302, 1297, 1293, 1289, 1285, 1280, 1276, 1272, 1267, 1263, 1259, 1254, 1250, 1245, 1240, 1236,
1231, 1227, 1222, 1217, 1213, 1208, 1203, 1198, 1194, 1189, 1184, 1179, 1174, 1170, 1165, 1160,
1155, 1150, 1145, 1140, 1135, 1131, 1126, 1121, 1116, 1111, 1106, 1101, 1096, 1091, 1086, 1081,
1076, 1071, 1066, 1061, 1057, 1052, 1047, 1042, 1037, 1032, 1027, 1022, 1017, 1012, 1007, 1003,
997, 993, 988, 983, 978, 974, 969, 963, 959, 955, 950, 945, 940, 936, 931, 925),
(1434, 1434, 1433, 1433, 1433, 1433, 1432, 1432, 1431, 1430, 1430, 1429, 1428, 1427, 1426, 1425,
1424, 1422, 1421, 1420, 1418, 1417, 1415, 1413, 1411, 1410, 1408, 1406, 1404, 1401, 1399, 1397,
1395, 1392, 1390, 1387, 1385, 1382, 1379, 1376, 1374, 1371, 1368, 1365, 1362, 1358, 1355, 1352,
1349, 1345, 1342, 1339, 1335, 1331, 1328, 1324, 1321, 1317, 1313, 1309, 1305, 1301, 1297, 1293,
1289, 1285, 1281, 1277, 1273, 1269, 1264, 1260, 1256, 1252, 1247, 1243, 1238, 1234, 1229, 1225,
1220, 1216, 1211, 1207, 1202, 1197, 1193, 1188, 1183, 1179, 1174, 1169, 1165, 1160, 1155, 1150,
1145, 1141, 1136, 1131, 1126, 1121, 1117, 1112, 1107, 1102, 1097, 1092, 1087, 1083, 1078, 1073,
1068, 1063, 1058, 1053, 1049, 1044, 1039, 1034, 1029, 1024, 1018, 1014, 1010, 1005, 1000, 995,
991, 986, 980, 976, 972, 967, 962, 957, 953, 948, 942, 939, 933, 929, 925, 920),
(1419, 1419, 1419, 1418, 1418, 1418, 1417, 1417, 1416, 1416, 1415, 1414, 1413, 1412, 1411, 1410,
1409, 1408, 1406, 1405, 1404, 1402, 1400, 1399, 1397, 1395, 1393, 1391, 1389, 1387, 1385, 1383,
1381, 1378, 1376, 1373, 1371, 1368, 1365, 1363, 1360, 1357, 1354, 1351, 1348, 1345, 1342, 1339,
1336, 1332, 1329, 1326, 1322, 1319, 1315, 1312, 1308, 1304, 1301, 1297, 1293, 1289, 1285, 1281,
1277, 1273, 1269, 1265, 1261, 1257, 1253, 1249, 1244, 1240, 1236, 1232, 1227, 1223, 1219, 1214,
1210, 1205, 1201, 1196, 1192, 1187, 1183, 1178, 1173, 1169, 1164, 1159, 1155, 1150, 1145, 1141,
1136, 1131, 1127, 1122, 1117, 1112, 1108, 1103, 1098, 1093, 1088, 1084, 1079, 1074, 1069, 1064,
1060, 1055, 1050, 1045, 1041, 1036, 1031, 1026, 1021, 1017, 1012, 1007, 1001, 997, 993, 988,
984, 979, 974, 969, 965, 959, 955, 950, 946, 941, 937, 932, 928, 923, 918, 914),
(1404, 1404, 1404, 1404, 1404, 1403, 1403, 1402, 1402, 1401, 1400, 1400, 1399, 1398, 1397, 1396,
1395, 1393, 1392, 1391, 1389, 1388, 1386, 1385, 1383, 1381, 1379, 1377, 1375, 1373, 1371, 1369,
1367, 1364, 1362, 1360, 1357, 1355, 1352, 1349, 1347, 1344, 1341, 1338, 1335, 1332, 1329, 1326,
1323, 1319, 1316, 1313, 1310, 1306, 1303, 1299, 1296, 1292, 1288, 1285, 1281, 1277, 1273, 1269,
1266, 1262, 1258, 1254, 1250, 1246, 1242, 1237, 1233, 1229, 1225, 1221, 1216, 1212, 1208, 1203,
1199, 1195, 1190, 1186, 1181, 1177, 1172, 1168, 1163, 1159, 1154, 1150, 1145, 1140, 1136, 1131,
1127, 1122, 1117, 1113, 1108, 1103, 1099, 1094, 1089, 1085, 1080, 1075, 1070, 1066, 1061, 1056,
1052, 1047, 1042, 1037, 1033, 1028, 1023, 1018, 1014, 1009, 1004, 1000, 995, 990, 986, 980,
976, 972, 967, 963, 958, 953, 949, 944, 940, 935, 929, 925, 921, 916, 912, 908),
(1390, 1390, 1390, 1389, 1389, 1389, 1388, 1388, 1387, 1387, 1386, 1385, 1385, 1384, 1383, 1382,
1380, 1379, 1378, 1377, 1375, 1374, 1372, 1371, 1369, 1367, 1365, 1363, 1362, 1360, 1357, 1355,
1353, 1351, 1349, 1346, 1344, 1341, 1339, 1336, 1333, 1331, 1328, 1325, 1322, 1319, 1316, 1313,
1310, 1307, 1304, 1300, 1297, 1294, 1290, 1287, 1283, 1280, 1276, 1273, 1269, 1265, 1261, 1258,
1254, 1250, 1246, 1242, 1238, 1234, 1230, 1226, 1222, 1218, 1214, 1210, 1206, 1201, 1197, 1193,
1189, 1184, 1180, 1176, 1171, 1167, 1162, 1158, 1153, 1149, 1145, 1140, 1135, 1131, 1126, 1122,
1117, 1113, 1108, 1104, 1099, 1094, 1090, 1085, 1081, 1076, 1071, 1067, 1062, 1057, 1053, 1048,
1043, 1039, 1034, 1030, 1025, 1020, 1016, 1010, 1006, 1001, 997, 992, 988, 983, 979, 974,
970, 965, 959, 956, 950, 946, 942, 938, 933, 929, 924, 920, 915, 911, 906, 902),
(1376, 1376, 1376, 1375, 1375, 1375, 1374, 1374, 1373, 1373, 1372, 1371, 1370, 1370, 1369, 1368,
1366, 1365, 1364, 1363, 1361, 1360, 1358, 1357, 1355, 1353, 1352, 1350, 1348, 1346, 1344, 1342,
1340, 1338, 1335, 1333, 1330, 1328, 1326, 1323, 1320, 1318, 1315, 1312, 1309, 1306, 1303, 1300,
1297, 1294, 1291, 1288, 1285, 1281, 1278, 1275, 1271, 1268, 1264, 1261, 1257, 1253, 1250, 1246,
1242, 1239, 1235, 1231, 1227, 1223, 1219, 1215, 1211, 1207, 1203, 1199, 1195, 1191, 1187, 1182,
1178, 1174, 1170, 1165, 1161, 1157, 1152, 1148, 1144, 1139, 1135, 1130, 1126, 1122, 1117, 1113,
1108, 1104, 1099, 1095, 1090, 1086, 1081, 1077, 1072, 1067, 1063, 1058, 1054, 1049, 1045, 1040,
1035, 1031, 1026, 1022, 1017, 1013, 1008, 1003, 999, 993, 990, 984, 980, 976, 972, 967,
963, 958, 954, 949, 945, 940, 936, 931, 927, 922, 918, 912, 909, 905, 899, 895),
(1362, 1362, 1362, 1361, 1361, 1361, 1360, 1360, 1359, 1359, 1358, 1357, 1357, 1356, 1355, 1354,
1353, 1352, 1350, 1349, 1348, 1346, 1345, 1343, 1342, 1340, 1338, 1336, 1335, 1333, 1331, 1329,
1327, 1324, 1322, 1320, 1317, 1315, 1313, 1310, 1307, 1305, 1302, 1299, 1297, 1294, 1291, 1288,
1285, 1282, 1279, 1276, 1273, 1269, 1266, 1263, 1259, 1256, 1252, 1249, 1245, 1242, 1238, 1235,
1231, 1227, 1224, 1220, 1216, 1212, 1208, 1204, 1200, 1196, 1192, 1188, 1184, 1180, 1176, 1172,
1168, 1164, 1160, 1155, 1151, 1147, 1143, 1138, 1134, 1130, 1125, 1121, 1117, 1112, 1108, 1104,
1099, 1095, 1090, 1086, 1081, 1077, 1072, 1068, 1064, 1059, 1055, 1050, 1046, 1041, 1037, 1032,
1028, 1023, 1018, 1014, 1010, 1005, 1001, 996, 992, 987, 983, 978, 974, 969, 965, 959,
956, 950, 946, 942, 938, 933, 929, 925, 920, 916, 912, 907, 903, 899, 894, 890),
(1348, 1348, 1348, 1348, 1347, 1347, 1347, 1346, 1346, 1345, 1345, 1344, 1343, 1342, 1341, 1340,
1339, 1338, 1337, 1336, 1334, 1333, 1331, 1330, 1328, 1327, 1325, 1323, 1321, 1320, 1318, 1316,
1313, 1311, 1309, 1307, 1305, 1302, 1300, 1297, 1295, 1292, 1290, 1287, 1284, 1281, 1279, 1276,
1273, 1270, 1267, 1264, 1261, 1257, 1254, 1251, 1248, 1244, 1241, 1237, 1234, 1230, 1227, 1223,
1220, 1216, 1212, 1209, 1205, 1201, 1197, 1194, 1190, 1186, 1182, 1178, 1174, 1170, 1166, 1162,
1158, 1154, 1150, 1145, 1141, 1137, 1133, 1129, 1125, 1120, 1116, 1112, 1107, 1103, 1099, 1094,
1090, 1086, 1081, 1077, 1073, 1068, 1064, 1060, 1055, 1051, 1046, 1042, 1037, 1033, 1029, 1024,
1020, 1014, 1010, 1006, 1001, 997, 993, 989, 984, 980, 975, 971, 967, 962, 958, 953,
949, 945, 940, 936, 931, 927, 923, 918, 914, 910, 905, 901, 897, 893, 888, 884),
(1334, 1334, 1334, 1334, 1334, 1334, 1333, 1333, 1332, 1332, 1331, 1330, 1330, 1329, 1328, 1327,
1326, 1325, 1324, 1322, 1321, 1320, 1318, 1317, 1315, 1314, 1312, 1310, 1308, 1307, 1305, 1303,
1301, 1299, 1296, 1294, 1292, 1290, 1287, 1285, 1282, 1280, 1277, 1275, 1272, 1269, 1266, 1264,
1261, 1258, 1255, 1252, 1249, 1246, 1242, 1239, 1236, 1233, 1229, 1226, 1223, 1219, 1216, 1212,
1209, 1205, 1202, 1198, 1194, 1190, 1187, 1183, 1179, 1175, 1172, 1168, 1164, 1160, 1156, 1152,
1148, 1144, 1140, 1136, 1132, 1128, 1123, 1119, 1115, 1111, 1107, 1103, 1098, 1094, 1090, 1086,
1081, 1077, 1073, 1068, 1064, 1060, 1055, 1051, 1047, 1042, 1038, 1034, 1029, 1025, 1021, 1016,
1012, 1008, 1003, 999, 993, 990, 986, 980, 976, 973, 967, 963, 959, 955, 950, 946,
942, 938, 933, 929, 925, 921, 916, 912, 908, 903, 899, 895, 891, 886, 882, 878),
(1321, 1321, 1321, 1321, 1321, 1320, 1320, 1320, 1319, 1318, 1318, 1317, 1316, 1316, 1315, 1314,
1313, 1312, 1310, 1309, 1308, 1307, 1305, 1304, 1302, 1301, 1299, 1297, 1296, 1294, 1292, 1290,
1288, 1286, 1284, 1282, 1279, 1277, 1275, 1272, 1270, 1268, 1265, 1262, 1260, 1257, 1254, 1252,
1249, 1246, 1243, 1240, 1237, 1234, 1231, 1228, 1225, 1221, 1218, 1215, 1211, 1208, 1205, 1201,
1198, 1194, 1191, 1187, 1184, 1180, 1176, 1173, 1169, 1165, 1161, 1157, 1154, 1150, 1146, 1142,
1138, 1134, 1130, 1126, 1122, 1118, 1114, 1110, 1106, 1102, 1098, 1093, 1089, 1085, 1081, 1077,
1073, 1068, 1064, 1060, 1056, 1051, 1047, 1043, 1039, 1034, 1030, 1026, 1021, 1017, 1013, 1009,
1004, 1000, 996, 991, 987, 983, 978, 974, 970, 966, 961, 957, 953, 948, 944, 940,
936, 931, 927, 923, 919, 914, 910, 906, 902, 897, 893, 889, 885, 881, 877, 872),
(1308, 1308, 1308, 1308, 1308, 1307, 1307, 1306, 1306, 1305, 1305, 1304, 1303, 1303, 1302, 1301,
1300, 1299, 1298, 1296, 1295, 1294, 1292, 1291, 1290, 1288, 1286, 1285, 1283, 1281, 1279, 1277,
1276, 1274, 1271, 1269, 1267, 1265, 1263, 1260, 1258, 1256, 1253, 1250, 1248, 1245, 1243, 1240,
1237, 1234, 1231, 1228, 1226, 1223, 1220, 1216, 1213, 1210, 1207, 1204, 1200, 1197, 1194, 1190,
1187, 1184, 1180, 1177, 1173, 1169, 1166, 1162, 1159, 1155, 1151, 1147, 1144, 1140, 1136, 1132,
1128, 1124, 1120, 1117, 1113, 1109, 1105, 1101, 1097, 1093, 1088, 1084, 1080, 1076, 1072, 1068,
1064, 1060, 1056, 1051, 1047, 1043, 1039, 1035, 1030, 1026, 1022, 1018, 1014, 1009, 1005, 1001,
997, 992, 988, 984, 980, 976, 971, 967, 963, 959, 954, 950, 946, 942, 937, 933,
929, 925, 921, 916, 912, 908, 903, 899, 895, 891, 886, 882, 878, 875, 871, 867),
(1295, 1295, 1295, 1295, 1295, 1294, 1294, 1294, 1293, 1293, 1292, 1291, 1291, 1290, 1289, 1288,
1287, 1286, 1285, 1284, 1282, 1281, 1280, 1278, 1277, 1275, 1274, 1272, 1271, 1269, 1267, 1265,
1263, 1261, 1259, 1257, 1255, 1253, 1251, 1248, 1246, 1244, 1241, 1239, 1236, 1234, 1231, 1228,
1226, 1223, 1220, 1217, 1214, 1211, 1208, 1205, 1202, 1199, 1196, 1193, 1190, 1186, 1183, 1180,
1176, 1173, 1170, 1166, 1163, 1159, 1156, 1152, 1148, 1145, 1141, 1137, 1134, 1130, 1126, 1122,
1119, 1115, 1111, 1107, 1103, 1099, 1095, 1091, 1087, 1084, 1080, 1076, 1072, 1067, 1063, 1059,
1055, 1051, 1047, 1043, 1039, 1035, 1031, 1027, 1022, 1018, 1014, 1010, 1006, 1001, 997, 993,
989, 984, 980, 976, 972, 967, 963, 959, 956, 952, 946, 942, 939, 935, 931, 927,
922, 918, 914, 910, 906, 902, 898, 894, 889, 885, 881, 877, 873, 869, 865, 861),
(1282, 1282, 1282, 1282, 1282, 1282, 1281, 1281, 1280, 1280, 1279, 1279, 1278, 1277, 1276, 1275,
1274, 1273, 1272, 1271, 1270, 1269, 1267, 1266, 1265, 1263, 1262, 1260, 1258, 1257, 1255, 1253,
1251, 1249, 1247, 1245, 1243, 1241, 1239, 1236, 1234, 1232, 1229, 1227, 1225, 1222, 1219, 1217,
1214, 1211, 1209, 1206, 1203, 1200, 1197, 1194, 1191, 1188, 1185, 1182, 1179, 1176, 1172, 1169,
1166, 1162, 1159, 1156, 1152, 1149, 1145, 1142, 1138, 1135, 1131, 1128, 1124, 1120, 1117, 1113,
1109, 1105, 1102, 1098, 1094, 1090, 1086, 1082, 1079, 1075, 1071, 1067, 1063, 1059, 1055, 1051,
1047, 1043, 1039, 1035, 1031, 1027, 1023, 1018, 1014, 1010, 1006, 1001, 997, 993, 990, 986,
982, 978, 974, 969, 965, 961, 957, 953, 949, 945, 941, 936, 932, 928, 924, 920,
916, 912, 908, 903, 899, 895, 892, 888, 882, 878, 875, 871, 867, 863, 859, 855),
(1270, 1270, 1270, 1270, 1269, 1269, 1269, 1268, 1268, 1267, 1267, 1266, 1265, 1265, 1264, 1263,
1262, 1261, 1260, 1259, 1258, 1256, 1255, 1254, 1252, 1251, 1249, 1248, 1246, 1245, 1243, 1241,
1239, 1237, 1235, 1233, 1231, 1229, 1227, 1225, 1223, 1220, 1218, 1216, 1213, 1211, 1208, 1205,
1203, 1200, 1197, 1195, 1192, 1189, 1186, 1183, 1180, 1177, 1174, 1171, 1168, 1165, 1162, 1159,
1155, 1152, 1149, 1146, 1142, 1139, 1135, 1132, 1128, 1125, 1121, 1118, 1114, 1111, 1107, 1103,
1100, 1096, 1092, 1089, 1085, 1081, 1077, 1073, 1070, 1066, 1062, 1058, 1054, 1050, 1046, 1042,
1038, 1035, 1031, 1027, 1023, 1018, 1014, 1010, 1007, 1003, 999, 995, 991, 987, 982, 978,
974, 970, 966, 962, 958, 954, 950, 946, 942, 938, 933, 929, 925, 922, 918, 914,
910, 906, 902, 898, 893, 889, 885, 881, 877, 874, 869, 865, 861, 858, 854, 850),
(1258, 1257, 1257, 1257, 1257, 1257, 1256, 1256, 1256, 1255, 1255, 1254, 1253, 1252, 1252, 1251,
1250, 1249, 1248, 1247, 1246, 1244, 1243, 1242, 1240, 1239, 1237, 1236, 1234, 1233, 1231, 1229,
1227, 1226, 1224, 1222, 1220, 1218, 1215, 1213, 1211, 1209, 1207, 1204, 1202, 1199, 1197, 1194,
1192, 1189, 1187, 1184, 1181, 1178, 1175, 1173, 1170, 1167, 1164, 1161, 1158, 1155, 1152, 1148,
1145, 1142, 1139, 1135, 1132, 1129, 1125, 1122, 1119, 1115, 1112, 1108, 1105, 1101, 1098, 1094,
1090, 1087, 1083, 1079, 1076, 1072, 1068, 1065, 1061, 1057, 1053, 1049, 1046, 1042, 1038, 1034,
1030, 1026, 1022, 1018, 1014, 1010, 1007, 1003, 999, 995, 991, 987, 983, 979, 975, 971,
967, 963, 959, 955, 950, 946, 942, 939, 935, 931, 927, 923, 919, 915, 911, 907,
903, 899, 895, 891, 886, 882, 878, 876, 872, 868, 864, 860, 856, 852, 848, 844),
(1245, 1245, 1245, 1245, 1245, 1245, 1244, 1244, 1243, 1243, 1242, 1242, 1241, 1240, 1240, 1239,
1238, 1237, 1236, 1235, 1234, 1232, 1231, 1230, 1229, 1227, 1226, 1224, 1223, 1221, 1219, 1218,
1216, 1214, 1212, 1210, 1208, 1206, 1204, 1202, 1200, 1198, 1195, 1193, 1191, 1188, 1186, 1183,
1181, 1178, 1176, 1173, 1170, 1168, 1165, 1162, 1159, 1156, 1153, 1150, 1147, 1144, 1141, 1138,
1135, 1132, 1129, 1126, 1122, 1119, 1116, 1112, 1109, 1106, 1102, 1099, 1095, 1092, 1088, 1085,
1081, 1078, 1074, 1070, 1067, 1063, 1060, 1056, 1052, 1048, 1045, 1041, 1037, 1033, 1030, 1026,
1022, 1018, 1014, 1010, 1007, 1003, 999, 995, 991, 987, 983, 979, 976, 972, 967, 963,
959, 956, 952, 948, 944, 940, 936, 932, 928, 924, 921, 916, 912, 909, 905, 901,
897, 893, 889, 885, 881, 877, 873, 869, 865, 861, 858, 854, 850, 846, 843, 839),
(1233, 1233, 1233, 1233, 1233, 1233, 1232, 1232, 1231, 1231, 1230, 1230, 1229, 1228, 1228, 1227,
1226, 1225, 1224, 1223, 1222, 1221, 1219, 1218, 1217, 1215, 1214, 1213, 1211, 1209, 1208, 1206,
1204, 1203, 1201, 1199, 1197, 1195, 1193, 1191, 1189, 1187, 1184, 1182, 1180, 1177, 1175, 1173,
1170, 1168, 1165, 1162, 1160, 1157, 1154, 1152, 1149, 1146, 1143, 1140, 1137, 1134, 1131, 1128,
1125, 1122, 1119, 1116, 1113, 1109, 1106, 1103, 1099, 1096, 1093, 1089, 1086, 1083, 1079, 1076,
1072, 1069, 1065, 1062, 1058, 1054, 1051, 1047, 1044, 1040, 1036, 1033, 1029, 1025, 1021, 1018,
1014, 1010, 1006, 1003, 999, 995, 991, 987, 984, 980, 976, 972, 967, 963, 959, 957,
953, 949, 945, 941, 937, 933, 929, 925, 922, 918, 914, 910, 906, 902, 898, 895,
891, 886, 882, 878, 875, 871, 868, 864, 860, 856, 852, 848, 844, 841, 837, 833),
(1222, 1221, 1221, 1221, 1221, 1221, 1220, 1220, 1220, 1219, 1219, 1218, 1217, 1217, 1216, 1215,
1214, 1213, 1212, 1211, 1210, 1209, 1208, 1207, 1205, 1204, 1203, 1201, 1200, 1198, 1196, 1195,
1193, 1191, 1190, 1188, 1186, 1184, 1182, 1180, 1178, 1176, 1173, 1171, 1169, 1167, 1164, 1162,
1159, 1157, 1154, 1152, 1149, 1147, 1144, 1141, 1138, 1136, 1133, 1130, 1127, 1124, 1121, 1118,
1115, 1112, 1109, 1106, 1103, 1100, 1097, 1093, 1090, 1087, 1084, 1080, 1077, 1073, 1070, 1067,
1063, 1060, 1056, 1053, 1049, 1046, 1042, 1039, 1035, 1031, 1028, 1024, 1021, 1017, 1013, 1010,
1006, 1001, 997, 995, 991, 987, 984, 980, 976, 972, 967, 965, 961, 957, 953, 949,
946, 942, 938, 933, 929, 927, 923, 919, 915, 911, 907, 903, 899, 895, 892, 888,
884, 881, 877, 873, 869, 865, 861, 858, 854, 850, 847, 843, 839, 835, 831, 827),
(1210, 1210, 1210, 1210, 1209, 1209, 1209, 1208, 1208, 1208, 1207, 1206, 1206, 1205, 1204, 1204,
1203, 1202, 1201, 1200, 1199, 1198, 1197, 1195, 1194, 1193, 1191, 1190, 1188, 1187, 1185, 1184,
1182, 1180, 1178, 1177, 1175, 1173, 1171, 1169, 1167, 1165, 1163, 1160, 1158, 1156, 1154, 1151,
1149, 1146, 1144, 1141, 1139, 1136, 1134, 1131, 1128, 1126, 1123, 1120, 1117, 1114, 1111, 1109,
1106, 1103, 1100, 1096, 1093, 1090, 1087, 1084, 1081, 1078, 1074, 1071, 1068, 1064, 1061, 1058,
1054, 1051, 1048, 1044, 1041, 1037, 1034, 1030, 1027, 1023, 1020, 1016, 1012, 1009, 1005, 1001,
997, 993, 991, 987, 983, 980, 976, 972, 969, 965, 961, 957, 954, 950, 946, 942,
939, 935, 931, 927, 924, 920, 916, 912, 909, 905, 901, 897, 893, 890, 886, 882,
878, 875, 871, 867, 863, 860, 856, 852, 848, 844, 841, 837, 834, 830, 826, 822),
(1198, 1198, 1198, 1198, 1198, 1198, 1197, 1197, 1197, 1196, 1196, 1195, 1194, 1194, 1193, 1192,
1191, 1190, 1190, 1189, 1188, 1186, 1185, 1184, 1183, 1182, 1180, 1179, 1177, 1176, 1174, 1173,
1171, 1169, 1168, 1166, 1164, 1162, 1160, 1158, 1156, 1154, 1152, 1150, 1148, 1145, 1143, 1141,
1139, 1136, 1134, 1131, 1129, 1126, 1124, 1121, 1118, 1116, 1113, 1110, 1107, 1105, 1102, 1099,
1096, 1093, 1090, 1087, 1084, 1081, 1078, 1075, 1072, 1068, 1065, 1062, 1059, 1056, 1052, 1049,
1046, 1042, 1039, 1036, 1032, 1029, 1025, 1022, 1018, 1014, 1010, 1008, 1004, 1001, 997, 993,
990, 987, 983, 979, 976, 972, 967, 965, 961, 958, 954, 950, 946, 942, 939, 935,
932, 928, 924, 921, 916, 912, 909, 906, 902, 898, 895, 891, 886, 882, 880, 876,
872, 869, 865, 861, 857, 854, 850, 846, 843, 839, 835, 831, 827, 824, 821, 817),
(1187, 1187, 1187, 1187, 1187, 1186, 1186, 1186, 1185, 1185, 1184, 1184, 1183, 1182, 1182, 1181,
1180, 1179, 1178, 1177, 1176, 1175, 1174, 1173, 1172, 1170, 1169, 1168, 1166, 1165, 1163, 1162,
1160, 1159, 1157, 1155, 1153, 1151, 1150, 1148, 1146, 1144, 1142, 1139, 1137, 1135, 1133, 1131,
1128, 1126, 1124, 1121, 1119, 1116, 1114, 1111, 1108, 1106, 1103, 1100, 1098, 1095, 1092, 1089,
1086, 1084, 1081, 1078, 1075, 1072, 1069, 1066, 1063, 1059, 1056, 1053, 1050, 1047, 1044, 1040,
1037, 1034, 1030, 1027, 1024, 1020, 1017, 1014, 1010, 1007, 1003, 1000, 996, 993, 989, 986,
982, 979, 975, 972, 967, 965, 961, 957, 954, 950, 946, 942, 939, 936, 932, 928,
925, 921, 918, 914, 910, 907, 903, 899, 895, 892, 888, 885, 881, 877, 874, 869,
865, 863, 859, 855, 852, 848, 844, 841, 837, 833, 830, 826, 823, 818, 814, 812),
(1176, 1176, 1176, 1176, 1175, 1175, 1175, 1175, 1174, 1174, 1173, 1173, 1172, 1171, 1171, 1170,
1169, 1168, 1167, 1166, 1165, 1164, 1163, 1162, 1161, 1160, 1158, 1157, 1156, 1154, 1153, 1151,
1149, 1148, 1146, 1144, 1143, 1141, 1139, 1137, 1135, 1133, 1131, 1129, 1127, 1125, 1123, 1120,
1118, 1116, 1114, 1111, 1109, 1106, 1104, 1101, 1099, 1096, 1093, 1091, 1088, 1085, 1083, 1080,
1077, 1074, 1071, 1068, 1066, 1063, 1060, 1057, 1054, 1051, 1047, 1044, 1041, 1038, 1035, 1032,
1028, 1025, 1022, 1018, 1014, 1012, 1009, 1005, 1001, 999, 995, 992, 989, 984, 982, 978,
975, 971, 967, 963, 961, 957, 954, 950, 946, 942, 940, 936, 932, 929, 925, 922,
918, 914, 911, 907, 903, 899, 895, 893, 889, 886, 882, 878, 875, 871, 868, 864,
860, 857, 852, 848, 846, 842, 839, 835, 831, 827, 824, 821, 817, 814, 810, 807),
(1165, 1165, 1165, 1165, 1164, 1164, 1164, 1164, 1163, 1163, 1162, 1162, 1161, 1160, 1160, 1159,
1158, 1157, 1157, 1156, 1155, 1154, 1152, 1151, 1150, 1149, 1148, 1146, 1145, 1144, 1142, 1141,
1139, 1137, 1136, 1134, 1132, 1131, 1129, 1127, 1125, 1123, 1121, 1119, 1117, 1115, 1113, 1110,
1108, 1106, 1104, 1101, 1099, 1097, 1094, 1092, 1089, 1087, 1084, 1081, 1079, 1076, 1073, 1071,
1068, 1065, 1062, 1059, 1056, 1054, 1051, 1048, 1045, 1042, 1039, 1036, 1033, 1029, 1026, 1023,
1020, 1017, 1014, 1010, 1007, 1004, 1001, 997, 993, 991, 987, 984, 980, 976, 974, 971,
967, 963, 959, 957, 953, 950, 946, 942, 939, 936, 932, 929, 925, 922, 918, 915,
911, 908, 903, 901, 897, 894, 890, 886, 882, 878, 876, 872, 869, 865, 861, 858,
854, 851, 847, 844, 840, 837, 833, 830, 826, 822, 818, 814, 812, 808, 805, 801),
(1154, 1154, 1154, 1154, 1154, 1153, 1153, 1153, 1152, 1152, 1151, 1151, 1150, 1150, 1149, 1148,
1148, 1147, 1146, 1145, 1144, 1143, 1142, 1141, 1140, 1138, 1137, 1136, 1134, 1133, 1132, 1130,
1129, 1127, 1125, 1124, 1122, 1120, 1118, 1117, 1115, 1113, 1111, 1109, 1107, 1105, 1103, 1101,
1098, 1096, 1094, 1092, 1089, 1087, 1084, 1082, 1080, 1077, 1075, 1072, 1069, 1067, 1064, 1061,
1059, 1056, 1053, 1050, 1048, 1045, 1042, 1039, 1036, 1033, 1030, 1027, 1024, 1021, 1018, 1014,
1012, 1009, 1005, 1001, 999, 996, 993, 989, 986, 983, 980, 976, 973, 970, 966, 963,
959, 956, 953, 950, 946, 942, 939, 936, 932, 929, 925, 922, 919, 915, 912, 908,
905, 901, 898, 894, 891, 886, 884, 880, 877, 873, 869, 865, 863, 859, 856, 852,
848, 844, 842, 838, 835, 831, 827, 824, 821, 817, 814, 810, 807, 803, 800, 796),
(1143, 1143, 1143, 1143, 1143, 1143, 1142, 1142, 1142, 1141, 1141, 1140, 1140, 1139, 1138, 1138,
1137, 1136, 1135, 1134, 1133, 1132, 1131, 1130, 1129, 1128, 1127, 1125, 1124, 1123, 1121, 1120,
1118, 1117, 1115, 1114, 1112, 1110, 1108, 1107, 1105, 1103, 1101, 1099, 1097, 1095, 1093, 1091,
1089, 1086, 1084, 1082, 1080, 1077, 1075, 1073, 1070, 1068, 1065, 1063, 1060, 1058, 1055, 1052,
1050, 1047, 1044, 1041, 1039, 1036, 1033, 1030, 1027, 1024, 1022, 1018, 1016, 1013, 1010, 1007,
1003, 1000, 997, 993, 991, 988, 984, 982, 978, 975, 972, 969, 965, 962, 959, 956,
952, 949, 946, 942, 939, 936, 932, 929, 925, 922, 919, 915, 912, 908, 905, 901,
898, 895, 891, 888, 884, 881, 877, 874, 869, 867, 864, 860, 857, 852, 850, 846,
843, 839, 835, 831, 829, 825, 822, 818, 814, 812, 808, 805, 801, 797, 795, 791),
(1133, 1133, 1133, 1132, 1132, 1132, 1132, 1132, 1131, 1131, 1130, 1130, 1129, 1129, 1128, 1127,
1126, 1126, 1125, 1124, 1123, 1122, 1121, 1120, 1119, 1118, 1116, 1115, 1114, 1113, 1111, 1110,
1108, 1107, 1105, 1104, 1102, 1100, 1098, 1097, 1095, 1093, 1091, 1089, 1087, 1085, 1083, 1081,
1079, 1077, 1075, 1073, 1070, 1068, 1066, 1063, 1061, 1059, 1056, 1054, 1051, 1049, 1046, 1043,
1041, 1038, 1035, 1033, 1030, 1027, 1024, 1022, 1018, 1016, 1013, 1010, 1007, 1004, 1001, 997,
995, 992, 989, 986, 983, 980, 976, 974, 971, 967, 963, 961, 958, 955, 950, 948,
945, 942, 938, 935, 932, 928, 925, 922, 918, 915, 912, 908, 905, 902, 898, 895,
892, 888, 885, 881, 878, 875, 871, 868, 864, 861, 857, 854, 851, 847, 844, 840,
837, 834, 830, 827, 823, 820, 817, 813, 810, 806, 803, 800, 796, 793, 789, 786),
(1122, 1122, 1122, 1122, 1122, 1122, 1121, 1121, 1121, 1120, 1120, 1119, 1119, 1118, 1118, 1117,
1116, 1115, 1115, 1114, 1113, 1112, 1111, 1110, 1109, 1107, 1106, 1105, 1104, 1102, 1101, 1100,
1098, 1097, 1095, 1094, 1092, 1090, 1089, 1087, 1085, 1083, 1082, 1080, 1078, 1076, 1074, 1072,
1070, 1068, 1065, 1063, 1061, 1059, 1056, 1054, 1052, 1049, 1047, 1045, 1042, 1040, 1037, 1035,
1032, 1029, 1027, 1024, 1021, 1018, 1016, 1013, 1010, 1008, 1005, 1001, 999, 996, 993, 990,
987, 984, 980, 978, 975, 972, 969, 966, 963, 959, 957, 954, 950, 946, 944, 941,
938, 933, 931, 928, 925, 921, 918, 915, 912, 908, 905, 902, 898, 895, 892, 888,
885, 882, 878, 875, 872, 868, 865, 861, 858, 855, 851, 848, 844, 841, 838, 835,
831, 827, 825, 821, 818, 814, 810, 808, 804, 801, 797, 793, 791, 788, 784, 781),
(1112, 1112, 1112, 1112, 1112, 1111, 1111, 1111, 1111, 1110, 1110, 1109, 1109, 1108, 1107, 1107,
1106, 1105, 1104, 1104, 1103, 1102, 1101, 1100, 1099, 1097, 1096, 1095, 1094, 1093, 1091, 1090,
1088, 1087, 1085, 1084, 1082, 1081, 1079, 1077, 1076, 1074, 1072, 1070, 1068, 1066, 1064, 1062,
1060, 1058, 1056, 1054, 1052, 1050, 1047, 1045, 1043, 1040, 1038, 1036, 1033, 1031, 1028, 1026,
1023, 1021, 1018, 1014, 1013, 1010, 1007, 1005, 1001, 999, 996, 993, 991, 988, 984, 982,
979, 976, 973, 970, 967, 963, 961, 958, 955, 952, 949, 946, 942, 940, 937, 933,
929, 927, 924, 921, 918, 915, 911, 908, 905, 902, 898, 895, 892, 889, 885, 882,
878, 875, 872, 869, 865, 861, 859, 856, 852, 848, 846, 842, 839, 835, 831, 829,
826, 822, 818, 816, 812, 809, 806, 801, 799, 796, 792, 789, 786, 783, 779, 776),
(1102, 1102, 1102, 1102, 1102, 1101, 1101, 1101, 1100, 1100, 1100, 1099, 1099, 1098, 1097, 1097,
1096, 1095, 1094, 1094, 1093, 1092, 1091, 1090, 1089, 1088, 1086, 1085, 1084, 1083, 1081, 1080,
1079, 1077, 1076, 1074, 1073, 1071, 1069, 1068, 1066, 1064, 1063, 1061, 1059, 1057, 1055, 1053,
1051, 1049, 1047, 1045, 1043, 1041, 1038, 1036, 1034, 1032, 1029, 1027, 1025, 1022, 1020, 1017,
1014, 1012, 1010, 1007, 1004, 1001, 999, 996, 993, 991, 988, 986, 983, 980, 976, 974,
971, 969, 966, 963, 959, 957, 954, 950, 948, 945, 942, 939, 936, 933, 929, 925,
923, 920, 916, 914, 911, 908, 903, 901, 898, 895, 892, 888, 885, 882, 878, 876,
872, 869, 865, 863, 859, 856, 852, 850, 846, 843, 840, 835, 833, 830, 827, 823,
820, 817, 813, 810, 807, 804, 800, 797, 793, 791, 787, 784, 781, 778, 774, 771),
(1092, 1092, 1092, 1092, 1092, 1091, 1091, 1091, 1090, 1090, 1090, 1089, 1089, 1088, 1087, 1087,
1086, 1085, 1085, 1084, 1083, 1082, 1081, 1080, 1079, 1078, 1077, 1076, 1074, 1073, 1072, 1070,
1069, 1068, 1066, 1065, 1063, 1062, 1060, 1058, 1057, 1055, 1053, 1051, 1050, 1048, 1046, 1044,
1042, 1040, 1038, 1036, 1034, 1032, 1029, 1027, 1025, 1023, 1021, 1018, 1016, 1013, 1010, 1009,
1006, 1004, 1001, 999, 996, 993, 991, 988, 986, 983, 980, 978, 975, 972, 969, 966,
963, 961, 958, 955, 952, 949, 946, 942, 940, 938, 935, 932, 929, 925, 922, 919,
916, 912, 910, 907, 903, 901, 898, 895, 891, 888, 885, 882, 878, 876, 872, 869,
865, 863, 860, 856, 852, 850, 847, 844, 840, 837, 834, 831, 827, 824, 821, 818,
814, 810, 808, 805, 801, 797, 795, 792, 789, 784, 782, 779, 776, 773, 769, 766),
(1082, 1082, 1082, 1082, 1082, 1081, 1081, 1081, 1081, 1080, 1080, 1079, 1079, 1078, 1078, 1077,
1076, 1076, 1075, 1074, 1073, 1072, 1071, 1070, 1069, 1068, 1067, 1066, 1065, 1064, 1062, 1061,
1060, 1058, 1057, 1055, 1054, 1052, 1051, 1049, 1047, 1046, 1044, 1042, 1041, 1039, 1037, 1035,
1033, 1031, 1029, 1027, 1025, 1023, 1021, 1018, 1016, 1014, 1012, 1010, 1007, 1005, 1003, 1000,
997, 995, 993, 990, 988, 984, 983, 980, 978, 975, 972, 970, 967, 963, 962, 959,
956, 953, 950, 948, 945, 942, 939, 936, 933, 929, 927, 924, 921, 918, 915, 912,
909, 906, 903, 899, 897, 894, 891, 888, 885, 882, 878, 876, 872, 869, 865, 863,
860, 857, 854, 850, 847, 844, 841, 838, 834, 831, 827, 825, 822, 818, 814, 812,
809, 806, 803, 799, 796, 793, 790, 787, 783, 780, 777, 774, 771, 768, 764, 761),
(1072, 1072, 1072, 1072, 1072, 1072, 1072, 1071, 1071, 1071, 1070, 1070, 1069, 1069, 1068, 1067,
1067, 1066, 1065, 1064, 1064, 1063, 1062, 1061, 1060, 1059, 1058, 1057, 1055, 1054, 1053, 1052,
1050, 1049, 1048, 1046, 1045, 1043, 1042, 1040, 1038, 1037, 1035, 1033, 1032, 1030, 1028, 1026,
1024, 1022, 1020, 1018, 1016, 1014, 1012, 1010, 1008, 1006, 1003, 1001, 999, 997, 993, 992,
990, 987, 984, 982, 980, 976, 975, 972, 970, 967, 963, 962, 959, 957, 954, 950,
948, 946, 942, 940, 937, 933, 932, 929, 925, 923, 920, 916, 914, 911, 908, 905,
902, 899, 897, 894, 891, 886, 884, 881, 878, 875, 872, 869, 865, 863, 860, 857,
854, 851, 847, 844, 841, 838, 835, 831, 829, 826, 822, 818, 816, 813, 810, 807,
804, 800, 797, 793, 791, 788, 784, 782, 778, 775, 772, 769, 766, 763, 760, 756),
(1063, 1063, 1063, 1063, 1062, 1062, 1062, 1062, 1061, 1061, 1061, 1060, 1060, 1059, 1059, 1058,
1057, 1057, 1056, 1055, 1054, 1053, 1052, 1051, 1050, 1049, 1048, 1047, 1046, 1045, 1044, 1042,
1041, 1040, 1038, 1037, 1036, 1034, 1033, 1031, 1029, 1028, 1026, 1024, 1023, 1021, 1018, 1017,
1014, 1013, 1012, 1010, 1008, 1006, 1003, 1001, 999, 997, 995, 993, 991, 988, 986, 984,
980, 979, 976, 974, 972, 969, 967, 963, 962, 959, 957, 954, 952, 949, 946, 944,
941, 938, 935, 933, 929, 927, 924, 922, 919, 916, 912, 910, 907, 903, 902, 899,
895, 893, 890, 886, 884, 881, 878, 875, 872, 869, 865, 863, 860, 857, 854, 851,
848, 844, 841, 838, 835, 831, 829, 826, 823, 820, 817, 814, 810, 807, 804, 801,
797, 795, 792, 789, 786, 783, 780, 776, 773, 770, 767, 764, 761, 758, 755, 752),
(1053, 1053, 1053, 1053, 1053, 1053, 1052, 1052, 1052, 1052, 1051, 1051, 1050, 1050, 1049, 1049,
1048, 1047, 1046, 1046, 1045, 1044, 1043, 1042, 1041, 1040, 1039, 1038, 1037, 1036, 1035, 1033,
1032, 1031, 1029, 1028, 1027, 1025, 1024, 1022, 1020, 1018, 1017, 1016, 1014, 1012, 1010, 1009,
1007, 1005, 1003, 1001, 999, 997, 995, 993, 991, 989, 987, 984, 982, 980, 978, 976,
973, 971, 969, 966, 963, 961, 959, 957, 954, 952, 949, 946, 944, 941, 939, 936,
933, 931, 928, 925, 923, 920, 916, 914, 912, 909, 906, 903, 899, 898, 895, 892,
889, 886, 882, 880, 877, 874, 871, 868, 865, 863, 860, 857, 854, 851, 848, 844,
842, 839, 835, 831, 829, 826, 823, 820, 817, 814, 810, 808, 805, 801, 799, 796,
793, 790, 787, 784, 781, 777, 774, 771, 768, 765, 762, 759, 756, 753, 750, 747),
(1044, 1044, 1044, 1044, 1044, 1043, 1043, 1043, 1043, 1042, 1042, 1041, 1041, 1040, 1040, 1039,
1039, 1038, 1037, 1036, 1036, 1035, 1034, 1033, 1032, 1031, 1030, 1029, 1028, 1027, 1026, 1024,
1023, 1022, 1020, 1018, 1018, 1016, 1014, 1013, 1012, 1010, 1009, 1007, 1005, 1004, 1001, 1000,
997, 996, 993, 993, 991, 989, 987, 984, 983, 980, 978, 976, 974, 972, 970, 967,
965, 963, 961, 958, 956, 954, 950, 949, 946, 944, 941, 939, 936, 933, 931, 929,
925, 923, 921, 918, 916, 912, 910, 907, 905, 902, 899, 895, 894, 891, 888, 885,
882, 878, 877, 874, 871, 868, 865, 861, 859, 856, 852, 850, 847, 844, 842, 839,
835, 833, 830, 827, 824, 821, 818, 814, 812, 809, 806, 803, 800, 797, 793, 790,
787, 784, 781, 778, 775, 772, 769, 766, 763, 760, 757, 754, 751, 748, 745, 742),
(1035, 1035, 1035, 1034, 1034, 1034, 1034, 1034, 1033, 1033, 1033, 1032, 1032, 1031, 1031, 1030,
1029, 1029, 1028, 1027, 1027, 1026, 1025, 1024, 1023, 1022, 1021, 1020, 1018, 1018, 1017, 1014,
1014, 1013, 1012, 1010, 1009, 1008, 1006, 1005, 1003, 1001, 1000, 997, 997, 995, 993, 992,
990, 988, 986, 984, 982, 980, 978, 976, 974, 972, 970, 967, 966, 963, 962, 959,
957, 955, 953, 950, 948, 946, 944, 941, 939, 936, 933, 931, 929, 925, 924, 921,
919, 916, 914, 911, 908, 906, 903, 899, 898, 895, 892, 890, 886, 884, 881, 878,
876, 873, 869, 867, 864, 861, 859, 856, 852, 850, 847, 844, 841, 838, 835, 833,
830, 827, 824, 821, 818, 814, 812, 809, 806, 803, 800, 797, 793, 791, 788, 784,
782, 779, 776, 773, 770, 767, 764, 761, 758, 755, 752, 749, 746, 743, 741, 738),
(1026, 1026, 1026, 1025, 1025, 1025, 1025, 1025, 1024, 1024, 1024, 1023, 1023, 1022, 1022, 1021,
1020, 1020, 1018, 1018, 1018, 1017, 1016, 1014, 1014, 1013, 1012, 1010, 1010, 1009, 1008, 1007,
1005, 1004, 1003, 1001, 1000, 999, 997, 996, 995, 993, 991, 990, 988, 987, 984, 983,
980, 980, 978, 976, 974, 972, 970, 967, 966, 963, 962, 959, 958, 956, 954, 952,
950, 946, 945, 942, 941, 938, 936, 933, 931, 929, 927, 924, 922, 919, 916, 914,
912, 909, 907, 903, 901, 899, 895, 894, 891, 888, 886, 882, 880, 877, 875, 872,
869, 865, 864, 861, 858, 855, 852, 850, 847, 844, 841, 838, 835, 831, 830, 827,
824, 821, 818, 814, 812, 809, 806, 803, 801, 797, 795, 792, 789, 786, 783, 780,
777, 774, 771, 768, 765, 762, 759, 756, 753, 751, 748, 745, 742, 739, 736, 733),
(1017, 1017, 1017, 1016, 1016, 1016, 1016, 1016, 1014, 1014, 1014, 1014, 1014, 1013, 1013, 1012,
1012, 1010, 1010, 1010, 1009, 1008, 1007, 1006, 1005, 1004, 1003, 1001, 1001, 1000, 999, 997,
997, 996, 993, 993, 992, 990, 989, 988, 986, 984, 983, 980, 980, 978, 976, 975,
973, 971, 970, 967, 966, 963, 962, 959, 958, 956, 954, 952, 950, 948, 946, 944,
942, 940, 938, 935, 933, 931, 929, 925, 924, 922, 919, 916, 914, 912, 910, 907,
905, 902, 899, 897, 894, 892, 889, 886, 884, 881, 878, 876, 874, 871, 868, 865,
863, 860, 857, 855, 852, 848, 846, 843, 841, 838, 835, 831, 829, 827, 824, 821,
818, 814, 812, 809, 807, 804, 801, 797, 795, 792, 789, 786, 783, 781, 778, 775,
772, 769, 766, 763, 760, 757, 754, 752, 749, 746, 743, 740, 737, 734, 731, 728),
(1008, 1008, 1008, 1008, 1007, 1007, 1007, 1007, 1007, 1006, 1006, 1005, 1005, 1004, 1004, 1003,
1003, 1001, 1001, 1001, 1000, 999, 997, 997, 997, 996, 995, 993, 993, 992, 991, 990,
988, 987, 986, 984, 983, 982, 980, 979, 978, 976, 975, 973, 972, 970, 967, 967,
965, 963, 962, 959, 958, 956, 954, 952, 950, 949, 946, 945, 942, 941, 939, 936,
933, 932, 929, 928, 925, 923, 921, 919, 916, 914, 912, 910, 907, 905, 902, 899,
898, 895, 893, 890, 888, 885, 882, 880, 877, 875, 872, 869, 867, 864, 861, 859,
856, 854, 851, 848, 846, 843, 840, 837, 835, 831, 829, 826, 823, 821, 818, 814,
812, 809, 807, 804, 801, 797, 795, 792, 790, 787, 784, 781, 778, 775, 772, 770,
767, 764, 761, 758, 755, 752, 750, 747, 744, 741, 738, 735, 732, 729, 727, 724)
);

constant EG_EG_INV_DR_SQ_LUT : calo_inv_dr_sq_lut_array := CALO_INV_DR_SQ_LUT;
constant EG_JET_INV_DR_SQ_LUT : calo_inv_dr_sq_lut_array := CALO_INV_DR_SQ_LUT;
constant EG_TAU_INV_DR_SQ_LUT : calo_inv_dr_sq_lut_array := CALO_INV_DR_SQ_LUT;
constant JET_JET_INV_DR_SQ_LUT : calo_inv_dr_sq_lut_array := CALO_INV_DR_SQ_LUT;
constant JET_TAU_INV_DR_SQ_LUT : calo_inv_dr_sq_lut_array := CALO_INV_DR_SQ_LUT;
constant TAU_TAU_INV_DR_SQ_LUT : calo_inv_dr_sq_lut_array := CALO_INV_DR_SQ_LUT;

end package;
