-- Description:
-- Package for LUTS with sfixed format values.

-- Version history:
-- HB 2020-03-14: first design

library ieee;
use ieee.std_logic_1164.all;
-- use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
-- use ieee.numeric_std.all;
use ieee.fixed_pkg.all;

-- use work.lhc_data_pkg.all;
-- use work.math_pkg.all;
use work.gtl_pkg.all;

package sfixed_luts_pkg is

type eg_pt_lut_sfixed_array is array (0 to 2**(D_S_I_EG_V2.et_high-D_S_I_EG_V2.et_low+1)-1) of sfixed(8 downto -20);
constant EG_PT_LUT_SFIXED : eg_pt_lut_sfixed_array := (
"00000000001001100110011001100", "00000000011001100110011001100", "00000000101001100110011001100", "00000000111001100110011001100", 
"00000001001001100110011001100", "00000001011001100110011001100", "00000001101001100110011001100", "00000001111001100110011001100", 
"00000010001001100110011001100", "00000010011001100110011001100", "00000010101001100110011001100", "00000010111001100110011001100", 
"00000011001001100110011001100", "00000011011001100110011001100", "00000011101001100110011001100", "00000011111001100110011001100", 
"00000100001001100110011001100", "00000100011001100110011001100", "00000100101001100110011001100", "00000100111001100110011001100", 
"00000101001001100110011001100", "00000101011001100110011001100", "00000101101001100110011001100", "00000101111001100110011001100", 
"00000110001001100110011001100", "00000110011001100110011001100", "00000110101001100110011001100", "00000110111001100110011001100", 
"00000111001001100110011001100", "00000111011001100110011001100", "00000111101001100110011001100", "00000111111001100110011001100", 
"00001000001001100110011001100", "00001000011001100110011001100", "00001000101001100110011001100", "00001000111001100110011001100", 
"00001001001001100110011001100", "00001001011001100110011001100", "00001001101001100110011001100", "00001001111001100110011001100", 
"00001010001001100110011001100", "00001010011001100110011001100", "00001010101001100110011001100", "00001010111001100110011001100", 
"00001011001001100110011001100", "00001011011001100110011001100", "00001011101001100110011001100", "00001011111001100110011001100", 
"00001100001001100110011001100", "00001100011001100110011001100", "00001100101001100110011001100", "00001100111001100110011001100", 
"00001101001001100110011001100", "00001101011001100110011001100", "00001101101001100110011001100", "00001101111001100110011001100", 
"00001110001001100110011001100", "00001110011001100110011001100", "00001110101001100110011001100", "00001110111001100110011001100", 
"00001111001001100110011001100", "00001111011001100110011001100", "00001111101001100110011001100", "00001111111001100110011001100", 
"00010000001001100110011001100", "00010000011001100110011001100", "00010000101001100110011001100", "00010000111001100110011001100", 
"00010001001001100110011001100", "00010001011001100110011001100", "00010001101001100110011001100", "00010001111001100110011001100", 
"00010010001001100110011001100", "00010010011001100110011001100", "00010010101001100110011001100", "00010010111001100110011001100", 
"00010011001001100110011001100", "00010011011001100110011001100", "00010011101001100110011001100", "00010011111001100110011001100", 
"00010100001001100110011001100", "00010100011001100110011001100", "00010100101001100110011001100", "00010100111001100110011001100", 
"00010101001001100110011001100", "00010101011001100110011001100", "00010101101001100110011001100", "00010101111001100110011001100", 
"00010110001001100110011001100", "00010110011001100110011001100", "00010110101001100110011001100", "00010110111001100110011001100", 
"00010111001001100110011001100", "00010111011001100110011001100", "00010111101001100110011001100", "00010111111001100110011001100", 
"00011000001001100110011001100", "00011000011001100110011001100", "00011000101001100110011001100", "00011000111001100110011001100", 
"00011001001001100110011001100", "00011001011001100110011001100", "00011001101001100110011001100", "00011001111001100110011001100", 
"00011010001001100110011001100", "00011010011001100110011001100", "00011010101001100110011001100", "00011010111001100110011001100", 
"00011011001001100110011001100", "00011011011001100110011001100", "00011011101001100110011001100", "00011011111001100110011001100", 
"00011100001001100110011001100", "00011100011001100110011001100", "00011100101001100110011001100", "00011100111001100110011001100", 
"00011101001001100110011001100", "00011101011001100110011001100", "00011101101001100110011001100", "00011101111001100110011001100", 
"00011110001001100110011001100", "00011110011001100110011001100", "00011110101001100110011001100", "00011110111001100110011001100", 
"00011111001001100110011001100", "00011111011001100110011001100", "00011111101001100110011001100", "00011111111001100110011001100", 
"00100000001001100110011001100", "00100000011001100110011001100", "00100000101001100110011001100", "00100000111001100110011001100", 
"00100001001001100110011001100", "00100001011001100110011001100", "00100001101001100110011001100", "00100001111001100110011001100", 
"00100010001001100110011001100", "00100010011001100110011001100", "00100010101001100110011001100", "00100010111001100110011001100", 
"00100011001001100110011001100", "00100011011001100110011001100", "00100011101001100110011001100", "00100011111001100110011001100", 
"00100100001001100110011001100", "00100100011001100110011001100", "00100100101001100110011001100", "00100100111001100110011001100", 
"00100101001001100110011001100", "00100101011001100110011001100", "00100101101001100110011001100", "00100101111001100110011001100", 
"00100110001001100110011001100", "00100110011001100110011001100", "00100110101001100110011001100", "00100110111001100110011001100", 
"00100111001001100110011001100", "00100111011001100110011001100", "00100111101001100110011001100", "00100111111001100110011001100", 
"00101000001001100110011001100", "00101000011001100110011001100", "00101000101001100110011001100", "00101000111001100110011001100", 
"00101001001001100110011001100", "00101001011001100110011001100", "00101001101001100110011001100", "00101001111001100110011001100", 
"00101010001001100110011001100", "00101010011001100110011001100", "00101010101001100110011001100", "00101010111001100110011001100", 
"00101011001001100110011001100", "00101011011001100110011001100", "00101011101001100110011001100", "00101011111001100110011001100", 
"00101100001001100110011001100", "00101100011001100110011001100", "00101100101001100110011001100", "00101100111001100110011001100", 
"00101101001001100110011001100", "00101101011001100110011001100", "00101101101001100110011001100", "00101101111001100110011001100", 
"00101110001001100110011001100", "00101110011001100110011001100", "00101110101001100110011001100", "00101110111001100110011001100", 
"00101111001001100110011001100", "00101111011001100110011001100", "00101111101001100110011001100", "00101111111001100110011001100", 
"00110000001001100110011001100", "00110000011001100110011001100", "00110000101001100110011001100", "00110000111001100110011001100", 
"00110001001001100110011001100", "00110001011001100110011001100", "00110001101001100110011001100", "00110001111001100110011001100", 
"00110010001001100110011001100", "00110010011001100110011001100", "00110010101001100110011001100", "00110010111001100110011001100", 
"00110011001001100110011001100", "00110011011001100110011001100", "00110011101001100110011001100", "00110011111001100110011001100", 
"00110100001001100110011001100", "00110100011001100110011001100", "00110100101001100110011001100", "00110100111001100110011001100", 
"00110101001001100110011001100", "00110101011001100110011001100", "00110101101001100110011001100", "00110101111001100110011001100", 
"00110110001001100110011001100", "00110110011001100110011001100", "00110110101001100110011001100", "00110110111001100110011001100", 
"00110111001001100110011001100", "00110111011001100110011001100", "00110111101001100110011001100", "00110111111001100110011001100", 
"00111000001001100110011001100", "00111000011001100110011001100", "00111000101001100110011001100", "00111000111001100110011001100", 
"00111001001001100110011001100", "00111001011001100110011001100", "00111001101001100110011001100", "00111001111001100110011001100", 
"00111010001001100110011001100", "00111010011001100110011001100", "00111010101001100110011001100", "00111010111001100110011001100", 
"00111011001001100110011001100", "00111011011001100110011001100", "00111011101001100110011001100", "00111011111001100110011001100", 
"00111100001001100110011001100", "00111100011001100110011001100", "00111100101001100110011001100", "00111100111001100110011001100", 
"00111101001001100110011001100", "00111101011001100110011001100", "00111101101001100110011001100", "00111101111001100110011001100", 
"00111110001001100110011001100", "00111110011001100110011001100", "00111110101001100110011001100", "00111110111001100110011001100", 
"00111111001001100110011001100", "00111111011001100110011001100", "00111111101001100110011001100", "00111111111001100110011001100", 
"01000000001001100110011001100", "01000000011001100110011001100", "01000000101001100110011001100", "01000000111001100110011001100", 
"01000001001001100110011001100", "01000001011001100110011001100", "01000001101001100110011001100", "01000001111001100110011001100", 
"01000010001001100110011001100", "01000010011001100110011001100", "01000010101001100110011001100", "01000010111001100110011001100", 
"01000011001001100110011001100", "01000011011001100110011001100", "01000011101001100110011001100", "01000011111001100110011001100", 
"01000100001001100110011001100", "01000100011001100110011001100", "01000100101001100110011001100", "01000100111001100110011001100", 
"01000101001001100110011001100", "01000101011001100110011001100", "01000101101001100110011001100", "01000101111001100110011001100", 
"01000110001001100110011001100", "01000110011001100110011001100", "01000110101001100110011001100", "01000110111001100110011001100", 
"01000111001001100110011001100", "01000111011001100110011001100", "01000111101001100110011001100", "01000111111001100110011001100", 
"01001000001001100110011001100", "01001000011001100110011001100", "01001000101001100110011001100", "01001000111001100110011001100", 
"01001001001001100110011001100", "01001001011001100110011001100", "01001001101001100110011001100", "01001001111001100110011001100", 
"01001010001001100110011001100", "01001010011001100110011001100", "01001010101001100110011001100", "01001010111001100110011001100", 
"01001011001001100110011001100", "01001011011001100110011001100", "01001011101001100110011001100", "01001011111001100110011001100", 
"01001100001001100110011001100", "01001100011001100110011001100", "01001100101001100110011001100", "01001100111001100110011001100", 
"01001101001001100110011001100", "01001101011001100110011001100", "01001101101001100110011001100", "01001101111001100110011001100", 
"01001110001001100110011001100", "01001110011001100110011001100", "01001110101001100110011001100", "01001110111001100110011001100", 
"01001111001001100110011001100", "01001111011001100110011001100", "01001111101001100110011001100", "01001111111001100110011001100", 
"01010000001001100110011001100", "01010000011001100110011001100", "01010000101001100110011001100", "01010000111001100110011001100", 
"01010001001001100110011001100", "01010001011001100110011001100", "01010001101001100110011001100", "01010001111001100110011001100", 
"01010010001001100110011001100", "01010010011001100110011001100", "01010010101001100110011001100", "01010010111001100110011001100", 
"01010011001001100110011001100", "01010011011001100110011001100", "01010011101001100110011001100", "01010011111001100110011001100", 
"01010100001001100110011001100", "01010100011001100110011001100", "01010100101001100110011001100", "01010100111001100110011001100", 
"01010101001001100110011001100", "01010101011001100110011001100", "01010101101001100110011001100", "01010101111001100110011001100", 
"01010110001001100110011001100", "01010110011001100110011001100", "01010110101001100110011001100", "01010110111001100110011001100", 
"01010111001001100110011001100", "01010111011001100110011001100", "01010111101001100110011001100", "01010111111001100110011001100", 
"01011000001001100110011001100", "01011000011001100110011001100", "01011000101001100110011001100", "01011000111001100110011001100", 
"01011001001001100110011001100", "01011001011001100110011001100", "01011001101001100110011001100", "01011001111001100110011001100", 
"01011010001001100110011001100", "01011010011001100110011001100", "01011010101001100110011001100", "01011010111001100110011001100", 
"01011011001001100110011001100", "01011011011001100110011001100", "01011011101001100110011001100", "01011011111001100110011001100", 
"01011100001001100110011001100", "01011100011001100110011001100", "01011100101001100110011001100", "01011100111001100110011001100", 
"01011101001001100110011001100", "01011101011001100110011001100", "01011101101001100110011001100", "01011101111001100110011001100", 
"01011110001001100110011001100", "01011110011001100110011001100", "01011110101001100110011001100", "01011110111001100110011001100", 
"01011111001001100110011001100", "01011111011001100110011001100", "01011111101001100110011001100", "01011111111001100110011001100", 
"01100000001001100110011001100", "01100000011001100110011001100", "01100000101001100110011001100", "01100000111001100110011001100", 
"01100001001001100110011001100", "01100001011001100110011001100", "01100001101001100110011001100", "01100001111001100110011001100", 
"01100010001001100110011001100", "01100010011001100110011001100", "01100010101001100110011001100", "01100010111001100110011001100", 
"01100011001001100110011001100", "01100011011001100110011001100", "01100011101001100110011001100", "01100011111001100110011001100", 
"01100100001001100110011001100", "01100100011001100110011001100", "01100100101001100110011001100", "01100100111001100110011001100", 
"01100101001001100110011001100", "01100101011001100110011001100", "01100101101001100110011001100", "01100101111001100110011001100", 
"01100110001001100110011001100", "01100110011001100110011001100", "01100110101001100110011001100", "01100110111001100110011001100", 
"01100111001001100110011001100", "01100111011001100110011001100", "01100111101001100110011001100", "01100111111001100110011001100", 
"01101000001001100110011001100", "01101000011001100110011001100", "01101000101001100110011001100", "01101000111001100110011001100", 
"01101001001001100110011001100", "01101001011001100110011001100", "01101001101001100110011001100", "01101001111001100110011001100", 
"01101010001001100110011001100", "01101010011001100110011001100", "01101010101001100110011001100", "01101010111001100110011001100", 
"01101011001001100110011001100", "01101011011001100110011001100", "01101011101001100110011001100", "01101011111001100110011001100", 
"01101100001001100110011001100", "01101100011001100110011001100", "01101100101001100110011001100", "01101100111001100110011001100", 
"01101101001001100110011001100", "01101101011001100110011001100", "01101101101001100110011001100", "01101101111001100110011001100", 
"01101110001001100110011001100", "01101110011001100110011001100", "01101110101001100110011001100", "01101110111001100110011001100", 
"01101111001001100110011001100", "01101111011001100110011001100", "01101111101001100110011001100", "01101111111001100110011001100", 
"01110000001001100110011001100", "01110000011001100110011001100", "01110000101001100110011001100", "01110000111001100110011001100", 
"01110001001001100110011001100", "01110001011001100110011001100", "01110001101001100110011001100", "01110001111001100110011001100", 
"01110010001001100110011001100", "01110010011001100110011001100", "01110010101001100110011001100", "01110010111001100110011001100", 
"01110011001001100110011001100", "01110011011001100110011001100", "01110011101001100110011001100", "01110011111001100110011001100", 
"01110100001001100110011001100", "01110100011001100110011001100", "01110100101001100110011001100", "01110100111001100110011001100", 
"01110101001001100110011001100", "01110101011001100110011001100", "01110101101001100110011001100", "01110101111001100110011001100", 
"01110110001001100110011001100", "01110110011001100110011001100", "01110110101001100110011001100", "01110110111001100110011001100", 
"01110111001001100110011001100", "01110111011001100110011001100", "01110111101001100110011001100", "01110111111001100110011001100", 
"01111000001001100110011001100", "01111000011001100110011001100", "01111000101001100110011001100", "01111000111001100110011001100", 
"01111001001001100110011001100", "01111001011001100110011001100", "01111001101001100110011001100", "01111001111001100110011001100", 
"01111010001001100110011001100", "01111010011001100110011001100", "01111010101001100110011001100", "01111010111001100110011001100", 
"01111011001001100110011001100", "01111011011001100110011001100", "01111011101001100110011001100", "01111011111001100110011001100", 
"01111100001001100110011001100", "01111100011001100110011001100", "01111100101001100110011001100", "01111100111001100110011001100", 
"01111101001001100110011001100", "01111101011001100110011001100", "01111101101001100110011001100", "01111101111001100110011001100", 
"01111110001001100110011001100", "01111110011001100110011001100", "01111110101001100110011001100", "01111110111001100110011001100", 
"01111111001001100110011001100", "01111111011001100110011001100", "01111111101001100110011001100", "01111111111001100110011001100"
);
type jet_pt_lut_sfixed_array is array (0 to 2**(D_S_I_JET_V2.et_high-D_S_I_JET_V2.et_low+1)-1) of sfixed(10 downto -20);
constant JET_PT_LUT_SFIXED : jet_pt_lut_sfixed_array := (
"0000000000001001100110011001100", "0000000000011001100110011001100", "0000000000101001100110011001100", "0000000000111001100110011001100", 
"0000000001001001100110011001100", "0000000001011001100110011001100", "0000000001101001100110011001100", "0000000001111001100110011001100", 
"0000000010001001100110011001100", "0000000010011001100110011001100", "0000000010101001100110011001100", "0000000010111001100110011001100", 
"0000000011001001100110011001100", "0000000011011001100110011001100", "0000000011101001100110011001100", "0000000011111001100110011001100", 
"0000000100001001100110011001100", "0000000100011001100110011001100", "0000000100101001100110011001100", "0000000100111001100110011001100", 
"0000000101001001100110011001100", "0000000101011001100110011001100", "0000000101101001100110011001100", "0000000101111001100110011001100", 
"0000000110001001100110011001100", "0000000110011001100110011001100", "0000000110101001100110011001100", "0000000110111001100110011001100", 
"0000000111001001100110011001100", "0000000111011001100110011001100", "0000000111101001100110011001100", "0000000111111001100110011001100", 
"0000001000001001100110011001100", "0000001000011001100110011001100", "0000001000101001100110011001100", "0000001000111001100110011001100", 
"0000001001001001100110011001100", "0000001001011001100110011001100", "0000001001101001100110011001100", "0000001001111001100110011001100", 
"0000001010001001100110011001100", "0000001010011001100110011001100", "0000001010101001100110011001100", "0000001010111001100110011001100", 
"0000001011001001100110011001100", "0000001011011001100110011001100", "0000001011101001100110011001100", "0000001011111001100110011001100", 
"0000001100001001100110011001100", "0000001100011001100110011001100", "0000001100101001100110011001100", "0000001100111001100110011001100", 
"0000001101001001100110011001100", "0000001101011001100110011001100", "0000001101101001100110011001100", "0000001101111001100110011001100", 
"0000001110001001100110011001100", "0000001110011001100110011001100", "0000001110101001100110011001100", "0000001110111001100110011001100", 
"0000001111001001100110011001100", "0000001111011001100110011001100", "0000001111101001100110011001100", "0000001111111001100110011001100", 
"0000010000001001100110011001100", "0000010000011001100110011001100", "0000010000101001100110011001100", "0000010000111001100110011001100", 
"0000010001001001100110011001100", "0000010001011001100110011001100", "0000010001101001100110011001100", "0000010001111001100110011001100", 
"0000010010001001100110011001100", "0000010010011001100110011001100", "0000010010101001100110011001100", "0000010010111001100110011001100", 
"0000010011001001100110011001100", "0000010011011001100110011001100", "0000010011101001100110011001100", "0000010011111001100110011001100", 
"0000010100001001100110011001100", "0000010100011001100110011001100", "0000010100101001100110011001100", "0000010100111001100110011001100", 
"0000010101001001100110011001100", "0000010101011001100110011001100", "0000010101101001100110011001100", "0000010101111001100110011001100", 
"0000010110001001100110011001100", "0000010110011001100110011001100", "0000010110101001100110011001100", "0000010110111001100110011001100", 
"0000010111001001100110011001100", "0000010111011001100110011001100", "0000010111101001100110011001100", "0000010111111001100110011001100", 
"0000011000001001100110011001100", "0000011000011001100110011001100", "0000011000101001100110011001100", "0000011000111001100110011001100", 
"0000011001001001100110011001100", "0000011001011001100110011001100", "0000011001101001100110011001100", "0000011001111001100110011001100", 
"0000011010001001100110011001100", "0000011010011001100110011001100", "0000011010101001100110011001100", "0000011010111001100110011001100", 
"0000011011001001100110011001100", "0000011011011001100110011001100", "0000011011101001100110011001100", "0000011011111001100110011001100", 
"0000011100001001100110011001100", "0000011100011001100110011001100", "0000011100101001100110011001100", "0000011100111001100110011001100", 
"0000011101001001100110011001100", "0000011101011001100110011001100", "0000011101101001100110011001100", "0000011101111001100110011001100", 
"0000011110001001100110011001100", "0000011110011001100110011001100", "0000011110101001100110011001100", "0000011110111001100110011001100", 
"0000011111001001100110011001100", "0000011111011001100110011001100", "0000011111101001100110011001100", "0000011111111001100110011001100", 
"0000100000001001100110011001100", "0000100000011001100110011001100", "0000100000101001100110011001100", "0000100000111001100110011001100", 
"0000100001001001100110011001100", "0000100001011001100110011001100", "0000100001101001100110011001100", "0000100001111001100110011001100", 
"0000100010001001100110011001100", "0000100010011001100110011001100", "0000100010101001100110011001100", "0000100010111001100110011001100", 
"0000100011001001100110011001100", "0000100011011001100110011001100", "0000100011101001100110011001100", "0000100011111001100110011001100", 
"0000100100001001100110011001100", "0000100100011001100110011001100", "0000100100101001100110011001100", "0000100100111001100110011001100", 
"0000100101001001100110011001100", "0000100101011001100110011001100", "0000100101101001100110011001100", "0000100101111001100110011001100", 
"0000100110001001100110011001100", "0000100110011001100110011001100", "0000100110101001100110011001100", "0000100110111001100110011001100", 
"0000100111001001100110011001100", "0000100111011001100110011001100", "0000100111101001100110011001100", "0000100111111001100110011001100", 
"0000101000001001100110011001100", "0000101000011001100110011001100", "0000101000101001100110011001100", "0000101000111001100110011001100", 
"0000101001001001100110011001100", "0000101001011001100110011001100", "0000101001101001100110011001100", "0000101001111001100110011001100", 
"0000101010001001100110011001100", "0000101010011001100110011001100", "0000101010101001100110011001100", "0000101010111001100110011001100", 
"0000101011001001100110011001100", "0000101011011001100110011001100", "0000101011101001100110011001100", "0000101011111001100110011001100", 
"0000101100001001100110011001100", "0000101100011001100110011001100", "0000101100101001100110011001100", "0000101100111001100110011001100", 
"0000101101001001100110011001100", "0000101101011001100110011001100", "0000101101101001100110011001100", "0000101101111001100110011001100", 
"0000101110001001100110011001100", "0000101110011001100110011001100", "0000101110101001100110011001100", "0000101110111001100110011001100", 
"0000101111001001100110011001100", "0000101111011001100110011001100", "0000101111101001100110011001100", "0000101111111001100110011001100", 
"0000110000001001100110011001100", "0000110000011001100110011001100", "0000110000101001100110011001100", "0000110000111001100110011001100", 
"0000110001001001100110011001100", "0000110001011001100110011001100", "0000110001101001100110011001100", "0000110001111001100110011001100", 
"0000110010001001100110011001100", "0000110010011001100110011001100", "0000110010101001100110011001100", "0000110010111001100110011001100", 
"0000110011001001100110011001100", "0000110011011001100110011001100", "0000110011101001100110011001100", "0000110011111001100110011001100", 
"0000110100001001100110011001100", "0000110100011001100110011001100", "0000110100101001100110011001100", "0000110100111001100110011001100", 
"0000110101001001100110011001100", "0000110101011001100110011001100", "0000110101101001100110011001100", "0000110101111001100110011001100", 
"0000110110001001100110011001100", "0000110110011001100110011001100", "0000110110101001100110011001100", "0000110110111001100110011001100", 
"0000110111001001100110011001100", "0000110111011001100110011001100", "0000110111101001100110011001100", "0000110111111001100110011001100", 
"0000111000001001100110011001100", "0000111000011001100110011001100", "0000111000101001100110011001100", "0000111000111001100110011001100", 
"0000111001001001100110011001100", "0000111001011001100110011001100", "0000111001101001100110011001100", "0000111001111001100110011001100", 
"0000111010001001100110011001100", "0000111010011001100110011001100", "0000111010101001100110011001100", "0000111010111001100110011001100", 
"0000111011001001100110011001100", "0000111011011001100110011001100", "0000111011101001100110011001100", "0000111011111001100110011001100", 
"0000111100001001100110011001100", "0000111100011001100110011001100", "0000111100101001100110011001100", "0000111100111001100110011001100", 
"0000111101001001100110011001100", "0000111101011001100110011001100", "0000111101101001100110011001100", "0000111101111001100110011001100", 
"0000111110001001100110011001100", "0000111110011001100110011001100", "0000111110101001100110011001100", "0000111110111001100110011001100", 
"0000111111001001100110011001100", "0000111111011001100110011001100", "0000111111101001100110011001100", "0000111111111001100110011001100", 
"0001000000001001100110011001100", "0001000000011001100110011001100", "0001000000101001100110011001100", "0001000000111001100110011001100", 
"0001000001001001100110011001100", "0001000001011001100110011001100", "0001000001101001100110011001100", "0001000001111001100110011001100", 
"0001000010001001100110011001100", "0001000010011001100110011001100", "0001000010101001100110011001100", "0001000010111001100110011001100", 
"0001000011001001100110011001100", "0001000011011001100110011001100", "0001000011101001100110011001100", "0001000011111001100110011001100", 
"0001000100001001100110011001100", "0001000100011001100110011001100", "0001000100101001100110011001100", "0001000100111001100110011001100", 
"0001000101001001100110011001100", "0001000101011001100110011001100", "0001000101101001100110011001100", "0001000101111001100110011001100", 
"0001000110001001100110011001100", "0001000110011001100110011001100", "0001000110101001100110011001100", "0001000110111001100110011001100", 
"0001000111001001100110011001100", "0001000111011001100110011001100", "0001000111101001100110011001100", "0001000111111001100110011001100", 
"0001001000001001100110011001100", "0001001000011001100110011001100", "0001001000101001100110011001100", "0001001000111001100110011001100", 
"0001001001001001100110011001100", "0001001001011001100110011001100", "0001001001101001100110011001100", "0001001001111001100110011001100", 
"0001001010001001100110011001100", "0001001010011001100110011001100", "0001001010101001100110011001100", "0001001010111001100110011001100", 
"0001001011001001100110011001100", "0001001011011001100110011001100", "0001001011101001100110011001100", "0001001011111001100110011001100", 
"0001001100001001100110011001100", "0001001100011001100110011001100", "0001001100101001100110011001100", "0001001100111001100110011001100", 
"0001001101001001100110011001100", "0001001101011001100110011001100", "0001001101101001100110011001100", "0001001101111001100110011001100", 
"0001001110001001100110011001100", "0001001110011001100110011001100", "0001001110101001100110011001100", "0001001110111001100110011001100", 
"0001001111001001100110011001100", "0001001111011001100110011001100", "0001001111101001100110011001100", "0001001111111001100110011001100", 
"0001010000001001100110011001100", "0001010000011001100110011001100", "0001010000101001100110011001100", "0001010000111001100110011001100", 
"0001010001001001100110011001100", "0001010001011001100110011001100", "0001010001101001100110011001100", "0001010001111001100110011001100", 
"0001010010001001100110011001100", "0001010010011001100110011001100", "0001010010101001100110011001100", "0001010010111001100110011001100", 
"0001010011001001100110011001100", "0001010011011001100110011001100", "0001010011101001100110011001100", "0001010011111001100110011001100", 
"0001010100001001100110011001100", "0001010100011001100110011001100", "0001010100101001100110011001100", "0001010100111001100110011001100", 
"0001010101001001100110011001100", "0001010101011001100110011001100", "0001010101101001100110011001100", "0001010101111001100110011001100", 
"0001010110001001100110011001100", "0001010110011001100110011001100", "0001010110101001100110011001100", "0001010110111001100110011001100", 
"0001010111001001100110011001100", "0001010111011001100110011001100", "0001010111101001100110011001100", "0001010111111001100110011001100", 
"0001011000001001100110011001100", "0001011000011001100110011001100", "0001011000101001100110011001100", "0001011000111001100110011001100", 
"0001011001001001100110011001100", "0001011001011001100110011001100", "0001011001101001100110011001100", "0001011001111001100110011001100", 
"0001011010001001100110011001100", "0001011010011001100110011001100", "0001011010101001100110011001100", "0001011010111001100110011001100", 
"0001011011001001100110011001100", "0001011011011001100110011001100", "0001011011101001100110011001100", "0001011011111001100110011001100", 
"0001011100001001100110011001100", "0001011100011001100110011001100", "0001011100101001100110011001100", "0001011100111001100110011001100", 
"0001011101001001100110011001100", "0001011101011001100110011001100", "0001011101101001100110011001100", "0001011101111001100110011001100", 
"0001011110001001100110011001100", "0001011110011001100110011001100", "0001011110101001100110011001100", "0001011110111001100110011001100", 
"0001011111001001100110011001100", "0001011111011001100110011001100", "0001011111101001100110011001100", "0001011111111001100110011001100", 
"0001100000001001100110011001100", "0001100000011001100110011001100", "0001100000101001100110011001100", "0001100000111001100110011001100", 
"0001100001001001100110011001100", "0001100001011001100110011001100", "0001100001101001100110011001100", "0001100001111001100110011001100", 
"0001100010001001100110011001100", "0001100010011001100110011001100", "0001100010101001100110011001100", "0001100010111001100110011001100", 
"0001100011001001100110011001100", "0001100011011001100110011001100", "0001100011101001100110011001100", "0001100011111001100110011001100", 
"0001100100001001100110011001100", "0001100100011001100110011001100", "0001100100101001100110011001100", "0001100100111001100110011001100", 
"0001100101001001100110011001100", "0001100101011001100110011001100", "0001100101101001100110011001100", "0001100101111001100110011001100", 
"0001100110001001100110011001100", "0001100110011001100110011001100", "0001100110101001100110011001100", "0001100110111001100110011001100", 
"0001100111001001100110011001100", "0001100111011001100110011001100", "0001100111101001100110011001100", "0001100111111001100110011001100", 
"0001101000001001100110011001100", "0001101000011001100110011001100", "0001101000101001100110011001100", "0001101000111001100110011001100", 
"0001101001001001100110011001100", "0001101001011001100110011001100", "0001101001101001100110011001100", "0001101001111001100110011001100", 
"0001101010001001100110011001100", "0001101010011001100110011001100", "0001101010101001100110011001100", "0001101010111001100110011001100", 
"0001101011001001100110011001100", "0001101011011001100110011001100", "0001101011101001100110011001100", "0001101011111001100110011001100", 
"0001101100001001100110011001100", "0001101100011001100110011001100", "0001101100101001100110011001100", "0001101100111001100110011001100", 
"0001101101001001100110011001100", "0001101101011001100110011001100", "0001101101101001100110011001100", "0001101101111001100110011001100", 
"0001101110001001100110011001100", "0001101110011001100110011001100", "0001101110101001100110011001100", "0001101110111001100110011001100", 
"0001101111001001100110011001100", "0001101111011001100110011001100", "0001101111101001100110011001100", "0001101111111001100110011001100", 
"0001110000001001100110011001100", "0001110000011001100110011001100", "0001110000101001100110011001100", "0001110000111001100110011001100", 
"0001110001001001100110011001100", "0001110001011001100110011001100", "0001110001101001100110011001100", "0001110001111001100110011001100", 
"0001110010001001100110011001100", "0001110010011001100110011001100", "0001110010101001100110011001100", "0001110010111001100110011001100", 
"0001110011001001100110011001100", "0001110011011001100110011001100", "0001110011101001100110011001100", "0001110011111001100110011001100", 
"0001110100001001100110011001100", "0001110100011001100110011001100", "0001110100101001100110011001100", "0001110100111001100110011001100", 
"0001110101001001100110011001100", "0001110101011001100110011001100", "0001110101101001100110011001100", "0001110101111001100110011001100", 
"0001110110001001100110011001100", "0001110110011001100110011001100", "0001110110101001100110011001100", "0001110110111001100110011001100", 
"0001110111001001100110011001100", "0001110111011001100110011001100", "0001110111101001100110011001100", "0001110111111001100110011001100", 
"0001111000001001100110011001100", "0001111000011001100110011001100", "0001111000101001100110011001100", "0001111000111001100110011001100", 
"0001111001001001100110011001100", "0001111001011001100110011001100", "0001111001101001100110011001100", "0001111001111001100110011001100", 
"0001111010001001100110011001100", "0001111010011001100110011001100", "0001111010101001100110011001100", "0001111010111001100110011001100", 
"0001111011001001100110011001100", "0001111011011001100110011001100", "0001111011101001100110011001100", "0001111011111001100110011001100", 
"0001111100001001100110011001100", "0001111100011001100110011001100", "0001111100101001100110011001100", "0001111100111001100110011001100", 
"0001111101001001100110011001100", "0001111101011001100110011001100", "0001111101101001100110011001100", "0001111101111001100110011001100", 
"0001111110001001100110011001100", "0001111110011001100110011001100", "0001111110101001100110011001100", "0001111110111001100110011001100", 
"0001111111001001100110011001100", "0001111111011001100110011001100", "0001111111101001100110011001100", "0001111111111001100110011001100", 
"0010000000001001100110011001100", "0010000000011001100110011001100", "0010000000101001100110011001100", "0010000000111001100110011001100", 
"0010000001001001100110011001100", "0010000001011001100110011001100", "0010000001101001100110011001100", "0010000001111001100110011001100", 
"0010000010001001100110011001100", "0010000010011001100110011001100", "0010000010101001100110011001100", "0010000010111001100110011001100", 
"0010000011001001100110011001100", "0010000011011001100110011001100", "0010000011101001100110011001100", "0010000011111001100110011001100", 
"0010000100001001100110011001100", "0010000100011001100110011001100", "0010000100101001100110011001100", "0010000100111001100110011001100", 
"0010000101001001100110011001100", "0010000101011001100110011001100", "0010000101101001100110011001100", "0010000101111001100110011001100", 
"0010000110001001100110011001100", "0010000110011001100110011001100", "0010000110101001100110011001100", "0010000110111001100110011001100", 
"0010000111001001100110011001100", "0010000111011001100110011001100", "0010000111101001100110011001100", "0010000111111001100110011001100", 
"0010001000001001100110011001100", "0010001000011001100110011001100", "0010001000101001100110011001100", "0010001000111001100110011001100", 
"0010001001001001100110011001100", "0010001001011001100110011001100", "0010001001101001100110011001100", "0010001001111001100110011001100", 
"0010001010001001100110011001100", "0010001010011001100110011001100", "0010001010101001100110011001100", "0010001010111001100110011001100", 
"0010001011001001100110011001100", "0010001011011001100110011001100", "0010001011101001100110011001100", "0010001011111001100110011001100", 
"0010001100001001100110011001100", "0010001100011001100110011001100", "0010001100101001100110011001100", "0010001100111001100110011001100", 
"0010001101001001100110011001100", "0010001101011001100110011001100", "0010001101101001100110011001100", "0010001101111001100110011001100", 
"0010001110001001100110011001100", "0010001110011001100110011001100", "0010001110101001100110011001100", "0010001110111001100110011001100", 
"0010001111001001100110011001100", "0010001111011001100110011001100", "0010001111101001100110011001100", "0010001111111001100110011001100", 
"0010010000001001100110011001100", "0010010000011001100110011001100", "0010010000101001100110011001100", "0010010000111001100110011001100", 
"0010010001001001100110011001100", "0010010001011001100110011001100", "0010010001101001100110011001100", "0010010001111001100110011001100", 
"0010010010001001100110011001100", "0010010010011001100110011001100", "0010010010101001100110011001100", "0010010010111001100110011001100", 
"0010010011001001100110011001100", "0010010011011001100110011001100", "0010010011101001100110011001100", "0010010011111001100110011001100", 
"0010010100001001100110011001100", "0010010100011001100110011001100", "0010010100101001100110011001100", "0010010100111001100110011001100", 
"0010010101001001100110011001100", "0010010101011001100110011001100", "0010010101101001100110011001100", "0010010101111001100110011001100", 
"0010010110001001100110011001100", "0010010110011001100110011001100", "0010010110101001100110011001100", "0010010110111001100110011001100", 
"0010010111001001100110011001100", "0010010111011001100110011001100", "0010010111101001100110011001100", "0010010111111001100110011001100", 
"0010011000001001100110011001100", "0010011000011001100110011001100", "0010011000101001100110011001100", "0010011000111001100110011001100", 
"0010011001001001100110011001100", "0010011001011001100110011001100", "0010011001101001100110011001100", "0010011001111001100110011001100", 
"0010011010001001100110011001100", "0010011010011001100110011001100", "0010011010101001100110011001100", "0010011010111001100110011001100", 
"0010011011001001100110011001100", "0010011011011001100110011001100", "0010011011101001100110011001100", "0010011011111001100110011001100", 
"0010011100001001100110011001100", "0010011100011001100110011001100", "0010011100101001100110011001100", "0010011100111001100110011001100", 
"0010011101001001100110011001100", "0010011101011001100110011001100", "0010011101101001100110011001100", "0010011101111001100110011001100", 
"0010011110001001100110011001100", "0010011110011001100110011001100", "0010011110101001100110011001100", "0010011110111001100110011001100", 
"0010011111001001100110011001100", "0010011111011001100110011001100", "0010011111101001100110011001100", "0010011111111001100110011001100", 
"0010100000001001100110011001100", "0010100000011001100110011001100", "0010100000101001100110011001100", "0010100000111001100110011001100", 
"0010100001001001100110011001100", "0010100001011001100110011001100", "0010100001101001100110011001100", "0010100001111001100110011001100", 
"0010100010001001100110011001100", "0010100010011001100110011001100", "0010100010101001100110011001100", "0010100010111001100110011001100", 
"0010100011001001100110011001100", "0010100011011001100110011001100", "0010100011101001100110011001100", "0010100011111001100110011001100", 
"0010100100001001100110011001100", "0010100100011001100110011001100", "0010100100101001100110011001100", "0010100100111001100110011001100", 
"0010100101001001100110011001100", "0010100101011001100110011001100", "0010100101101001100110011001100", "0010100101111001100110011001100", 
"0010100110001001100110011001100", "0010100110011001100110011001100", "0010100110101001100110011001100", "0010100110111001100110011001100", 
"0010100111001001100110011001100", "0010100111011001100110011001100", "0010100111101001100110011001100", "0010100111111001100110011001100", 
"0010101000001001100110011001100", "0010101000011001100110011001100", "0010101000101001100110011001100", "0010101000111001100110011001100", 
"0010101001001001100110011001100", "0010101001011001100110011001100", "0010101001101001100110011001100", "0010101001111001100110011001100", 
"0010101010001001100110011001100", "0010101010011001100110011001100", "0010101010101001100110011001100", "0010101010111001100110011001100", 
"0010101011001001100110011001100", "0010101011011001100110011001100", "0010101011101001100110011001100", "0010101011111001100110011001100", 
"0010101100001001100110011001100", "0010101100011001100110011001100", "0010101100101001100110011001100", "0010101100111001100110011001100", 
"0010101101001001100110011001100", "0010101101011001100110011001100", "0010101101101001100110011001100", "0010101101111001100110011001100", 
"0010101110001001100110011001100", "0010101110011001100110011001100", "0010101110101001100110011001100", "0010101110111001100110011001100", 
"0010101111001001100110011001100", "0010101111011001100110011001100", "0010101111101001100110011001100", "0010101111111001100110011001100", 
"0010110000001001100110011001100", "0010110000011001100110011001100", "0010110000101001100110011001100", "0010110000111001100110011001100", 
"0010110001001001100110011001100", "0010110001011001100110011001100", "0010110001101001100110011001100", "0010110001111001100110011001100", 
"0010110010001001100110011001100", "0010110010011001100110011001100", "0010110010101001100110011001100", "0010110010111001100110011001100", 
"0010110011001001100110011001100", "0010110011011001100110011001100", "0010110011101001100110011001100", "0010110011111001100110011001100", 
"0010110100001001100110011001100", "0010110100011001100110011001100", "0010110100101001100110011001100", "0010110100111001100110011001100", 
"0010110101001001100110011001100", "0010110101011001100110011001100", "0010110101101001100110011001100", "0010110101111001100110011001100", 
"0010110110001001100110011001100", "0010110110011001100110011001100", "0010110110101001100110011001100", "0010110110111001100110011001100", 
"0010110111001001100110011001100", "0010110111011001100110011001100", "0010110111101001100110011001100", "0010110111111001100110011001100", 
"0010111000001001100110011001100", "0010111000011001100110011001100", "0010111000101001100110011001100", "0010111000111001100110011001100", 
"0010111001001001100110011001100", "0010111001011001100110011001100", "0010111001101001100110011001100", "0010111001111001100110011001100", 
"0010111010001001100110011001100", "0010111010011001100110011001100", "0010111010101001100110011001100", "0010111010111001100110011001100", 
"0010111011001001100110011001100", "0010111011011001100110011001100", "0010111011101001100110011001100", "0010111011111001100110011001100", 
"0010111100001001100110011001100", "0010111100011001100110011001100", "0010111100101001100110011001100", "0010111100111001100110011001100", 
"0010111101001001100110011001100", "0010111101011001100110011001100", "0010111101101001100110011001100", "0010111101111001100110011001100", 
"0010111110001001100110011001100", "0010111110011001100110011001100", "0010111110101001100110011001100", "0010111110111001100110011001100", 
"0010111111001001100110011001100", "0010111111011001100110011001100", "0010111111101001100110011001100", "0010111111111001100110011001100", 
"0011000000001001100110011001100", "0011000000011001100110011001100", "0011000000101001100110011001100", "0011000000111001100110011001100", 
"0011000001001001100110011001100", "0011000001011001100110011001100", "0011000001101001100110011001100", "0011000001111001100110011001100", 
"0011000010001001100110011001100", "0011000010011001100110011001100", "0011000010101001100110011001100", "0011000010111001100110011001100", 
"0011000011001001100110011001100", "0011000011011001100110011001100", "0011000011101001100110011001100", "0011000011111001100110011001100", 
"0011000100001001100110011001100", "0011000100011001100110011001100", "0011000100101001100110011001100", "0011000100111001100110011001100", 
"0011000101001001100110011001100", "0011000101011001100110011001100", "0011000101101001100110011001100", "0011000101111001100110011001100", 
"0011000110001001100110011001100", "0011000110011001100110011001100", "0011000110101001100110011001100", "0011000110111001100110011001100", 
"0011000111001001100110011001100", "0011000111011001100110011001100", "0011000111101001100110011001100", "0011000111111001100110011001100", 
"0011001000001001100110011001100", "0011001000011001100110011001100", "0011001000101001100110011001100", "0011001000111001100110011001100", 
"0011001001001001100110011001100", "0011001001011001100110011001100", "0011001001101001100110011001100", "0011001001111001100110011001100", 
"0011001010001001100110011001100", "0011001010011001100110011001100", "0011001010101001100110011001100", "0011001010111001100110011001100", 
"0011001011001001100110011001100", "0011001011011001100110011001100", "0011001011101001100110011001100", "0011001011111001100110011001100", 
"0011001100001001100110011001100", "0011001100011001100110011001100", "0011001100101001100110011001100", "0011001100111001100110011001100", 
"0011001101001001100110011001100", "0011001101011001100110011001100", "0011001101101001100110011001100", "0011001101111001100110011001100", 
"0011001110001001100110011001100", "0011001110011001100110011001100", "0011001110101001100110011001100", "0011001110111001100110011001100", 
"0011001111001001100110011001100", "0011001111011001100110011001100", "0011001111101001100110011001100", "0011001111111001100110011001100", 
"0011010000001001100110011001100", "0011010000011001100110011001100", "0011010000101001100110011001100", "0011010000111001100110011001100", 
"0011010001001001100110011001100", "0011010001011001100110011001100", "0011010001101001100110011001100", "0011010001111001100110011001100", 
"0011010010001001100110011001100", "0011010010011001100110011001100", "0011010010101001100110011001100", "0011010010111001100110011001100", 
"0011010011001001100110011001100", "0011010011011001100110011001100", "0011010011101001100110011001100", "0011010011111001100110011001100", 
"0011010100001001100110011001100", "0011010100011001100110011001100", "0011010100101001100110011001100", "0011010100111001100110011001100", 
"0011010101001001100110011001100", "0011010101011001100110011001100", "0011010101101001100110011001100", "0011010101111001100110011001100", 
"0011010110001001100110011001100", "0011010110011001100110011001100", "0011010110101001100110011001100", "0011010110111001100110011001100", 
"0011010111001001100110011001100", "0011010111011001100110011001100", "0011010111101001100110011001100", "0011010111111001100110011001100", 
"0011011000001001100110011001100", "0011011000011001100110011001100", "0011011000101001100110011001100", "0011011000111001100110011001100", 
"0011011001001001100110011001100", "0011011001011001100110011001100", "0011011001101001100110011001100", "0011011001111001100110011001100", 
"0011011010001001100110011001100", "0011011010011001100110011001100", "0011011010101001100110011001100", "0011011010111001100110011001100", 
"0011011011001001100110011001100", "0011011011011001100110011001100", "0011011011101001100110011001100", "0011011011111001100110011001100", 
"0011011100001001100110011001100", "0011011100011001100110011001100", "0011011100101001100110011001100", "0011011100111001100110011001100", 
"0011011101001001100110011001100", "0011011101011001100110011001100", "0011011101101001100110011001100", "0011011101111001100110011001100", 
"0011011110001001100110011001100", "0011011110011001100110011001100", "0011011110101001100110011001100", "0011011110111001100110011001100", 
"0011011111001001100110011001100", "0011011111011001100110011001100", "0011011111101001100110011001100", "0011011111111001100110011001100", 
"0011100000001001100110011001100", "0011100000011001100110011001100", "0011100000101001100110011001100", "0011100000111001100110011001100", 
"0011100001001001100110011001100", "0011100001011001100110011001100", "0011100001101001100110011001100", "0011100001111001100110011001100", 
"0011100010001001100110011001100", "0011100010011001100110011001100", "0011100010101001100110011001100", "0011100010111001100110011001100", 
"0011100011001001100110011001100", "0011100011011001100110011001100", "0011100011101001100110011001100", "0011100011111001100110011001100", 
"0011100100001001100110011001100", "0011100100011001100110011001100", "0011100100101001100110011001100", "0011100100111001100110011001100", 
"0011100101001001100110011001100", "0011100101011001100110011001100", "0011100101101001100110011001100", "0011100101111001100110011001100", 
"0011100110001001100110011001100", "0011100110011001100110011001100", "0011100110101001100110011001100", "0011100110111001100110011001100", 
"0011100111001001100110011001100", "0011100111011001100110011001100", "0011100111101001100110011001100", "0011100111111001100110011001100", 
"0011101000001001100110011001100", "0011101000011001100110011001100", "0011101000101001100110011001100", "0011101000111001100110011001100", 
"0011101001001001100110011001100", "0011101001011001100110011001100", "0011101001101001100110011001100", "0011101001111001100110011001100", 
"0011101010001001100110011001100", "0011101010011001100110011001100", "0011101010101001100110011001100", "0011101010111001100110011001100", 
"0011101011001001100110011001100", "0011101011011001100110011001100", "0011101011101001100110011001100", "0011101011111001100110011001100", 
"0011101100001001100110011001100", "0011101100011001100110011001100", "0011101100101001100110011001100", "0011101100111001100110011001100", 
"0011101101001001100110011001100", "0011101101011001100110011001100", "0011101101101001100110011001100", "0011101101111001100110011001100", 
"0011101110001001100110011001100", "0011101110011001100110011001100", "0011101110101001100110011001100", "0011101110111001100110011001100", 
"0011101111001001100110011001100", "0011101111011001100110011001100", "0011101111101001100110011001100", "0011101111111001100110011001100", 
"0011110000001001100110011001100", "0011110000011001100110011001100", "0011110000101001100110011001100", "0011110000111001100110011001100", 
"0011110001001001100110011001100", "0011110001011001100110011001100", "0011110001101001100110011001100", "0011110001111001100110011001100", 
"0011110010001001100110011001100", "0011110010011001100110011001100", "0011110010101001100110011001100", "0011110010111001100110011001100", 
"0011110011001001100110011001100", "0011110011011001100110011001100", "0011110011101001100110011001100", "0011110011111001100110011001100", 
"0011110100001001100110011001100", "0011110100011001100110011001100", "0011110100101001100110011001100", "0011110100111001100110011001100", 
"0011110101001001100110011001100", "0011110101011001100110011001100", "0011110101101001100110011001100", "0011110101111001100110011001100", 
"0011110110001001100110011001100", "0011110110011001100110011001100", "0011110110101001100110011001100", "0011110110111001100110011001100", 
"0011110111001001100110011001100", "0011110111011001100110011001100", "0011110111101001100110011001100", "0011110111111001100110011001100", 
"0011111000001001100110011001100", "0011111000011001100110011001100", "0011111000101001100110011001100", "0011111000111001100110011001100", 
"0011111001001001100110011001100", "0011111001011001100110011001100", "0011111001101001100110011001100", "0011111001111001100110011001100", 
"0011111010001001100110011001100", "0011111010011001100110011001100", "0011111010101001100110011001100", "0011111010111001100110011001100", 
"0011111011001001100110011001100", "0011111011011001100110011001100", "0011111011101001100110011001100", "0011111011111001100110011001100", 
"0011111100001001100110011001100", "0011111100011001100110011001100", "0011111100101001100110011001100", "0011111100111001100110011001100", 
"0011111101001001100110011001100", "0011111101011001100110011001100", "0011111101101001100110011001100", "0011111101111001100110011001100", 
"0011111110001001100110011001100", "0011111110011001100110011001100", "0011111110101001100110011001100", "0011111110111001100110011001100", 
"0011111111001001100110011001100", "0011111111011001100110011001100", "0011111111101001100110011001100", "0011111111111001100110011001100", 
"0100000000001001100110011001100", "0100000000011001100110011001100", "0100000000101001100110011001100", "0100000000111001100110011001100", 
"0100000001001001100110011001100", "0100000001011001100110011001100", "0100000001101001100110011001100", "0100000001111001100110011001100", 
"0100000010001001100110011001100", "0100000010011001100110011001100", "0100000010101001100110011001100", "0100000010111001100110011001100", 
"0100000011001001100110011001100", "0100000011011001100110011001100", "0100000011101001100110011001100", "0100000011111001100110011001100", 
"0100000100001001100110011001100", "0100000100011001100110011001100", "0100000100101001100110011001100", "0100000100111001100110011001100", 
"0100000101001001100110011001100", "0100000101011001100110011001100", "0100000101101001100110011001100", "0100000101111001100110011001100", 
"0100000110001001100110011001100", "0100000110011001100110011001100", "0100000110101001100110011001100", "0100000110111001100110011001100", 
"0100000111001001100110011001100", "0100000111011001100110011001100", "0100000111101001100110011001100", "0100000111111001100110011001100", 
"0100001000001001100110011001100", "0100001000011001100110011001100", "0100001000101001100110011001100", "0100001000111001100110011001100", 
"0100001001001001100110011001100", "0100001001011001100110011001100", "0100001001101001100110011001100", "0100001001111001100110011001100", 
"0100001010001001100110011001100", "0100001010011001100110011001100", "0100001010101001100110011001100", "0100001010111001100110011001100", 
"0100001011001001100110011001100", "0100001011011001100110011001100", "0100001011101001100110011001100", "0100001011111001100110011001100", 
"0100001100001001100110011001100", "0100001100011001100110011001100", "0100001100101001100110011001100", "0100001100111001100110011001100", 
"0100001101001001100110011001100", "0100001101011001100110011001100", "0100001101101001100110011001100", "0100001101111001100110011001100", 
"0100001110001001100110011001100", "0100001110011001100110011001100", "0100001110101001100110011001100", "0100001110111001100110011001100", 
"0100001111001001100110011001100", "0100001111011001100110011001100", "0100001111101001100110011001100", "0100001111111001100110011001100", 
"0100010000001001100110011001100", "0100010000011001100110011001100", "0100010000101001100110011001100", "0100010000111001100110011001100", 
"0100010001001001100110011001100", "0100010001011001100110011001100", "0100010001101001100110011001100", "0100010001111001100110011001100", 
"0100010010001001100110011001100", "0100010010011001100110011001100", "0100010010101001100110011001100", "0100010010111001100110011001100", 
"0100010011001001100110011001100", "0100010011011001100110011001100", "0100010011101001100110011001100", "0100010011111001100110011001100", 
"0100010100001001100110011001100", "0100010100011001100110011001100", "0100010100101001100110011001100", "0100010100111001100110011001100", 
"0100010101001001100110011001100", "0100010101011001100110011001100", "0100010101101001100110011001100", "0100010101111001100110011001100", 
"0100010110001001100110011001100", "0100010110011001100110011001100", "0100010110101001100110011001100", "0100010110111001100110011001100", 
"0100010111001001100110011001100", "0100010111011001100110011001100", "0100010111101001100110011001100", "0100010111111001100110011001100", 
"0100011000001001100110011001100", "0100011000011001100110011001100", "0100011000101001100110011001100", "0100011000111001100110011001100", 
"0100011001001001100110011001100", "0100011001011001100110011001100", "0100011001101001100110011001100", "0100011001111001100110011001100", 
"0100011010001001100110011001100", "0100011010011001100110011001100", "0100011010101001100110011001100", "0100011010111001100110011001100", 
"0100011011001001100110011001100", "0100011011011001100110011001100", "0100011011101001100110011001100", "0100011011111001100110011001100", 
"0100011100001001100110011001100", "0100011100011001100110011001100", "0100011100101001100110011001100", "0100011100111001100110011001100", 
"0100011101001001100110011001100", "0100011101011001100110011001100", "0100011101101001100110011001100", "0100011101111001100110011001100", 
"0100011110001001100110011001100", "0100011110011001100110011001100", "0100011110101001100110011001100", "0100011110111001100110011001100", 
"0100011111001001100110011001100", "0100011111011001100110011001100", "0100011111101001100110011001100", "0100011111111001100110011001100", 
"0100100000001001100110011001100", "0100100000011001100110011001100", "0100100000101001100110011001100", "0100100000111001100110011001100", 
"0100100001001001100110011001100", "0100100001011001100110011001100", "0100100001101001100110011001100", "0100100001111001100110011001100", 
"0100100010001001100110011001100", "0100100010011001100110011001100", "0100100010101001100110011001100", "0100100010111001100110011001100", 
"0100100011001001100110011001100", "0100100011011001100110011001100", "0100100011101001100110011001100", "0100100011111001100110011001100", 
"0100100100001001100110011001100", "0100100100011001100110011001100", "0100100100101001100110011001100", "0100100100111001100110011001100", 
"0100100101001001100110011001100", "0100100101011001100110011001100", "0100100101101001100110011001100", "0100100101111001100110011001100", 
"0100100110001001100110011001100", "0100100110011001100110011001100", "0100100110101001100110011001100", "0100100110111001100110011001100", 
"0100100111001001100110011001100", "0100100111011001100110011001100", "0100100111101001100110011001100", "0100100111111001100110011001100", 
"0100101000001001100110011001100", "0100101000011001100110011001100", "0100101000101001100110011001100", "0100101000111001100110011001100", 
"0100101001001001100110011001100", "0100101001011001100110011001100", "0100101001101001100110011001100", "0100101001111001100110011001100", 
"0100101010001001100110011001100", "0100101010011001100110011001100", "0100101010101001100110011001100", "0100101010111001100110011001100", 
"0100101011001001100110011001100", "0100101011011001100110011001100", "0100101011101001100110011001100", "0100101011111001100110011001100", 
"0100101100001001100110011001100", "0100101100011001100110011001100", "0100101100101001100110011001100", "0100101100111001100110011001100", 
"0100101101001001100110011001100", "0100101101011001100110011001100", "0100101101101001100110011001100", "0100101101111001100110011001100", 
"0100101110001001100110011001100", "0100101110011001100110011001100", "0100101110101001100110011001100", "0100101110111001100110011001100", 
"0100101111001001100110011001100", "0100101111011001100110011001100", "0100101111101001100110011001100", "0100101111111001100110011001100", 
"0100110000001001100110011001100", "0100110000011001100110011001100", "0100110000101001100110011001100", "0100110000111001100110011001100", 
"0100110001001001100110011001100", "0100110001011001100110011001100", "0100110001101001100110011001100", "0100110001111001100110011001100", 
"0100110010001001100110011001100", "0100110010011001100110011001100", "0100110010101001100110011001100", "0100110010111001100110011001100", 
"0100110011001001100110011001100", "0100110011011001100110011001100", "0100110011101001100110011001100", "0100110011111001100110011001100", 
"0100110100001001100110011001100", "0100110100011001100110011001100", "0100110100101001100110011001100", "0100110100111001100110011001100", 
"0100110101001001100110011001100", "0100110101011001100110011001100", "0100110101101001100110011001100", "0100110101111001100110011001100", 
"0100110110001001100110011001100", "0100110110011001100110011001100", "0100110110101001100110011001100", "0100110110111001100110011001100", 
"0100110111001001100110011001100", "0100110111011001100110011001100", "0100110111101001100110011001100", "0100110111111001100110011001100", 
"0100111000001001100110011001100", "0100111000011001100110011001100", "0100111000101001100110011001100", "0100111000111001100110011001100", 
"0100111001001001100110011001100", "0100111001011001100110011001100", "0100111001101001100110011001100", "0100111001111001100110011001100", 
"0100111010001001100110011001100", "0100111010011001100110011001100", "0100111010101001100110011001100", "0100111010111001100110011001100", 
"0100111011001001100110011001100", "0100111011011001100110011001100", "0100111011101001100110011001100", "0100111011111001100110011001100", 
"0100111100001001100110011001100", "0100111100011001100110011001100", "0100111100101001100110011001100", "0100111100111001100110011001100", 
"0100111101001001100110011001100", "0100111101011001100110011001100", "0100111101101001100110011001100", "0100111101111001100110011001100", 
"0100111110001001100110011001100", "0100111110011001100110011001100", "0100111110101001100110011001100", "0100111110111001100110011001100", 
"0100111111001001100110011001100", "0100111111011001100110011001100", "0100111111101001100110011001100", "0100111111111001100110011001100", 
"0101000000001001100110011001100", "0101000000011001100110011001100", "0101000000101001100110011001100", "0101000000111001100110011001100", 
"0101000001001001100110011001100", "0101000001011001100110011001100", "0101000001101001100110011001100", "0101000001111001100110011001100", 
"0101000010001001100110011001100", "0101000010011001100110011001100", "0101000010101001100110011001100", "0101000010111001100110011001100", 
"0101000011001001100110011001100", "0101000011011001100110011001100", "0101000011101001100110011001100", "0101000011111001100110011001100", 
"0101000100001001100110011001100", "0101000100011001100110011001100", "0101000100101001100110011001100", "0101000100111001100110011001100", 
"0101000101001001100110011001100", "0101000101011001100110011001100", "0101000101101001100110011001100", "0101000101111001100110011001100", 
"0101000110001001100110011001100", "0101000110011001100110011001100", "0101000110101001100110011001100", "0101000110111001100110011001100", 
"0101000111001001100110011001100", "0101000111011001100110011001100", "0101000111101001100110011001100", "0101000111111001100110011001100", 
"0101001000001001100110011001100", "0101001000011001100110011001100", "0101001000101001100110011001100", "0101001000111001100110011001100", 
"0101001001001001100110011001100", "0101001001011001100110011001100", "0101001001101001100110011001100", "0101001001111001100110011001100", 
"0101001010001001100110011001100", "0101001010011001100110011001100", "0101001010101001100110011001100", "0101001010111001100110011001100", 
"0101001011001001100110011001100", "0101001011011001100110011001100", "0101001011101001100110011001100", "0101001011111001100110011001100", 
"0101001100001001100110011001100", "0101001100011001100110011001100", "0101001100101001100110011001100", "0101001100111001100110011001100", 
"0101001101001001100110011001100", "0101001101011001100110011001100", "0101001101101001100110011001100", "0101001101111001100110011001100", 
"0101001110001001100110011001100", "0101001110011001100110011001100", "0101001110101001100110011001100", "0101001110111001100110011001100", 
"0101001111001001100110011001100", "0101001111011001100110011001100", "0101001111101001100110011001100", "0101001111111001100110011001100", 
"0101010000001001100110011001100", "0101010000011001100110011001100", "0101010000101001100110011001100", "0101010000111001100110011001100", 
"0101010001001001100110011001100", "0101010001011001100110011001100", "0101010001101001100110011001100", "0101010001111001100110011001100", 
"0101010010001001100110011001100", "0101010010011001100110011001100", "0101010010101001100110011001100", "0101010010111001100110011001100", 
"0101010011001001100110011001100", "0101010011011001100110011001100", "0101010011101001100110011001100", "0101010011111001100110011001100", 
"0101010100001001100110011001100", "0101010100011001100110011001100", "0101010100101001100110011001100", "0101010100111001100110011001100", 
"0101010101001001100110011001100", "0101010101011001100110011001100", "0101010101101001100110011001100", "0101010101111001100110011001100", 
"0101010110001001100110011001100", "0101010110011001100110011001100", "0101010110101001100110011001100", "0101010110111001100110011001100", 
"0101010111001001100110011001100", "0101010111011001100110011001100", "0101010111101001100110011001100", "0101010111111001100110011001100", 
"0101011000001001100110011001100", "0101011000011001100110011001100", "0101011000101001100110011001100", "0101011000111001100110011001100", 
"0101011001001001100110011001100", "0101011001011001100110011001100", "0101011001101001100110011001100", "0101011001111001100110011001100", 
"0101011010001001100110011001100", "0101011010011001100110011001100", "0101011010101001100110011001100", "0101011010111001100110011001100", 
"0101011011001001100110011001100", "0101011011011001100110011001100", "0101011011101001100110011001100", "0101011011111001100110011001100", 
"0101011100001001100110011001100", "0101011100011001100110011001100", "0101011100101001100110011001100", "0101011100111001100110011001100", 
"0101011101001001100110011001100", "0101011101011001100110011001100", "0101011101101001100110011001100", "0101011101111001100110011001100", 
"0101011110001001100110011001100", "0101011110011001100110011001100", "0101011110101001100110011001100", "0101011110111001100110011001100", 
"0101011111001001100110011001100", "0101011111011001100110011001100", "0101011111101001100110011001100", "0101011111111001100110011001100", 
"0101100000001001100110011001100", "0101100000011001100110011001100", "0101100000101001100110011001100", "0101100000111001100110011001100", 
"0101100001001001100110011001100", "0101100001011001100110011001100", "0101100001101001100110011001100", "0101100001111001100110011001100", 
"0101100010001001100110011001100", "0101100010011001100110011001100", "0101100010101001100110011001100", "0101100010111001100110011001100", 
"0101100011001001100110011001100", "0101100011011001100110011001100", "0101100011101001100110011001100", "0101100011111001100110011001100", 
"0101100100001001100110011001100", "0101100100011001100110011001100", "0101100100101001100110011001100", "0101100100111001100110011001100", 
"0101100101001001100110011001100", "0101100101011001100110011001100", "0101100101101001100110011001100", "0101100101111001100110011001100", 
"0101100110001001100110011001100", "0101100110011001100110011001100", "0101100110101001100110011001100", "0101100110111001100110011001100", 
"0101100111001001100110011001100", "0101100111011001100110011001100", "0101100111101001100110011001100", "0101100111111001100110011001100", 
"0101101000001001100110011001100", "0101101000011001100110011001100", "0101101000101001100110011001100", "0101101000111001100110011001100", 
"0101101001001001100110011001100", "0101101001011001100110011001100", "0101101001101001100110011001100", "0101101001111001100110011001100", 
"0101101010001001100110011001100", "0101101010011001100110011001100", "0101101010101001100110011001100", "0101101010111001100110011001100", 
"0101101011001001100110011001100", "0101101011011001100110011001100", "0101101011101001100110011001100", "0101101011111001100110011001100", 
"0101101100001001100110011001100", "0101101100011001100110011001100", "0101101100101001100110011001100", "0101101100111001100110011001100", 
"0101101101001001100110011001100", "0101101101011001100110011001100", "0101101101101001100110011001100", "0101101101111001100110011001100", 
"0101101110001001100110011001100", "0101101110011001100110011001100", "0101101110101001100110011001100", "0101101110111001100110011001100", 
"0101101111001001100110011001100", "0101101111011001100110011001100", "0101101111101001100110011001100", "0101101111111001100110011001100", 
"0101110000001001100110011001100", "0101110000011001100110011001100", "0101110000101001100110011001100", "0101110000111001100110011001100", 
"0101110001001001100110011001100", "0101110001011001100110011001100", "0101110001101001100110011001100", "0101110001111001100110011001100", 
"0101110010001001100110011001100", "0101110010011001100110011001100", "0101110010101001100110011001100", "0101110010111001100110011001100", 
"0101110011001001100110011001100", "0101110011011001100110011001100", "0101110011101001100110011001100", "0101110011111001100110011001100", 
"0101110100001001100110011001100", "0101110100011001100110011001100", "0101110100101001100110011001100", "0101110100111001100110011001100", 
"0101110101001001100110011001100", "0101110101011001100110011001100", "0101110101101001100110011001100", "0101110101111001100110011001100", 
"0101110110001001100110011001100", "0101110110011001100110011001100", "0101110110101001100110011001100", "0101110110111001100110011001100", 
"0101110111001001100110011001100", "0101110111011001100110011001100", "0101110111101001100110011001100", "0101110111111001100110011001100", 
"0101111000001001100110011001100", "0101111000011001100110011001100", "0101111000101001100110011001100", "0101111000111001100110011001100", 
"0101111001001001100110011001100", "0101111001011001100110011001100", "0101111001101001100110011001100", "0101111001111001100110011001100", 
"0101111010001001100110011001100", "0101111010011001100110011001100", "0101111010101001100110011001100", "0101111010111001100110011001100", 
"0101111011001001100110011001100", "0101111011011001100110011001100", "0101111011101001100110011001100", "0101111011111001100110011001100", 
"0101111100001001100110011001100", "0101111100011001100110011001100", "0101111100101001100110011001100", "0101111100111001100110011001100", 
"0101111101001001100110011001100", "0101111101011001100110011001100", "0101111101101001100110011001100", "0101111101111001100110011001100", 
"0101111110001001100110011001100", "0101111110011001100110011001100", "0101111110101001100110011001100", "0101111110111001100110011001100", 
"0101111111001001100110011001100", "0101111111011001100110011001100", "0101111111101001100110011001100", "0101111111111001100110011001100", 
"0110000000001001100110011001100", "0110000000011001100110011001100", "0110000000101001100110011001100", "0110000000111001100110011001100", 
"0110000001001001100110011001100", "0110000001011001100110011001100", "0110000001101001100110011001100", "0110000001111001100110011001100", 
"0110000010001001100110011001100", "0110000010011001100110011001100", "0110000010101001100110011001100", "0110000010111001100110011001100", 
"0110000011001001100110011001100", "0110000011011001100110011001100", "0110000011101001100110011001100", "0110000011111001100110011001100", 
"0110000100001001100110011001100", "0110000100011001100110011001100", "0110000100101001100110011001100", "0110000100111001100110011001100", 
"0110000101001001100110011001100", "0110000101011001100110011001100", "0110000101101001100110011001100", "0110000101111001100110011001100", 
"0110000110001001100110011001100", "0110000110011001100110011001100", "0110000110101001100110011001100", "0110000110111001100110011001100", 
"0110000111001001100110011001100", "0110000111011001100110011001100", "0110000111101001100110011001100", "0110000111111001100110011001100", 
"0110001000001001100110011001100", "0110001000011001100110011001100", "0110001000101001100110011001100", "0110001000111001100110011001100", 
"0110001001001001100110011001100", "0110001001011001100110011001100", "0110001001101001100110011001100", "0110001001111001100110011001100", 
"0110001010001001100110011001100", "0110001010011001100110011001100", "0110001010101001100110011001100", "0110001010111001100110011001100", 
"0110001011001001100110011001100", "0110001011011001100110011001100", "0110001011101001100110011001100", "0110001011111001100110011001100", 
"0110001100001001100110011001100", "0110001100011001100110011001100", "0110001100101001100110011001100", "0110001100111001100110011001100", 
"0110001101001001100110011001100", "0110001101011001100110011001100", "0110001101101001100110011001100", "0110001101111001100110011001100", 
"0110001110001001100110011001100", "0110001110011001100110011001100", "0110001110101001100110011001100", "0110001110111001100110011001100", 
"0110001111001001100110011001100", "0110001111011001100110011001100", "0110001111101001100110011001100", "0110001111111001100110011001100", 
"0110010000001001100110011001100", "0110010000011001100110011001100", "0110010000101001100110011001100", "0110010000111001100110011001100", 
"0110010001001001100110011001100", "0110010001011001100110011001100", "0110010001101001100110011001100", "0110010001111001100110011001100", 
"0110010010001001100110011001100", "0110010010011001100110011001100", "0110010010101001100110011001100", "0110010010111001100110011001100", 
"0110010011001001100110011001100", "0110010011011001100110011001100", "0110010011101001100110011001100", "0110010011111001100110011001100", 
"0110010100001001100110011001100", "0110010100011001100110011001100", "0110010100101001100110011001100", "0110010100111001100110011001100", 
"0110010101001001100110011001100", "0110010101011001100110011001100", "0110010101101001100110011001100", "0110010101111001100110011001100", 
"0110010110001001100110011001100", "0110010110011001100110011001100", "0110010110101001100110011001100", "0110010110111001100110011001100", 
"0110010111001001100110011001100", "0110010111011001100110011001100", "0110010111101001100110011001100", "0110010111111001100110011001100", 
"0110011000001001100110011001100", "0110011000011001100110011001100", "0110011000101001100110011001100", "0110011000111001100110011001100", 
"0110011001001001100110011001100", "0110011001011001100110011001100", "0110011001101001100110011001100", "0110011001111001100110011001100", 
"0110011010001001100110011001100", "0110011010011001100110011001100", "0110011010101001100110011001100", "0110011010111001100110011001100", 
"0110011011001001100110011001100", "0110011011011001100110011001100", "0110011011101001100110011001100", "0110011011111001100110011001100", 
"0110011100001001100110011001100", "0110011100011001100110011001100", "0110011100101001100110011001100", "0110011100111001100110011001100", 
"0110011101001001100110011001100", "0110011101011001100110011001100", "0110011101101001100110011001100", "0110011101111001100110011001100", 
"0110011110001001100110011001100", "0110011110011001100110011001100", "0110011110101001100110011001100", "0110011110111001100110011001100", 
"0110011111001001100110011001100", "0110011111011001100110011001100", "0110011111101001100110011001100", "0110011111111001100110011001100", 
"0110100000001001100110011001100", "0110100000011001100110011001100", "0110100000101001100110011001100", "0110100000111001100110011001100", 
"0110100001001001100110011001100", "0110100001011001100110011001100", "0110100001101001100110011001100", "0110100001111001100110011001100", 
"0110100010001001100110011001100", "0110100010011001100110011001100", "0110100010101001100110011001100", "0110100010111001100110011001100", 
"0110100011001001100110011001100", "0110100011011001100110011001100", "0110100011101001100110011001100", "0110100011111001100110011001100", 
"0110100100001001100110011001100", "0110100100011001100110011001100", "0110100100101001100110011001100", "0110100100111001100110011001100", 
"0110100101001001100110011001100", "0110100101011001100110011001100", "0110100101101001100110011001100", "0110100101111001100110011001100", 
"0110100110001001100110011001100", "0110100110011001100110011001100", "0110100110101001100110011001100", "0110100110111001100110011001100", 
"0110100111001001100110011001100", "0110100111011001100110011001100", "0110100111101001100110011001100", "0110100111111001100110011001100", 
"0110101000001001100110011001100", "0110101000011001100110011001100", "0110101000101001100110011001100", "0110101000111001100110011001100", 
"0110101001001001100110011001100", "0110101001011001100110011001100", "0110101001101001100110011001100", "0110101001111001100110011001100", 
"0110101010001001100110011001100", "0110101010011001100110011001100", "0110101010101001100110011001100", "0110101010111001100110011001100", 
"0110101011001001100110011001100", "0110101011011001100110011001100", "0110101011101001100110011001100", "0110101011111001100110011001100", 
"0110101100001001100110011001100", "0110101100011001100110011001100", "0110101100101001100110011001100", "0110101100111001100110011001100", 
"0110101101001001100110011001100", "0110101101011001100110011001100", "0110101101101001100110011001100", "0110101101111001100110011001100", 
"0110101110001001100110011001100", "0110101110011001100110011001100", "0110101110101001100110011001100", "0110101110111001100110011001100", 
"0110101111001001100110011001100", "0110101111011001100110011001100", "0110101111101001100110011001100", "0110101111111001100110011001100", 
"0110110000001001100110011001100", "0110110000011001100110011001100", "0110110000101001100110011001100", "0110110000111001100110011001100", 
"0110110001001001100110011001100", "0110110001011001100110011001100", "0110110001101001100110011001100", "0110110001111001100110011001100", 
"0110110010001001100110011001100", "0110110010011001100110011001100", "0110110010101001100110011001100", "0110110010111001100110011001100", 
"0110110011001001100110011001100", "0110110011011001100110011001100", "0110110011101001100110011001100", "0110110011111001100110011001100", 
"0110110100001001100110011001100", "0110110100011001100110011001100", "0110110100101001100110011001100", "0110110100111001100110011001100", 
"0110110101001001100110011001100", "0110110101011001100110011001100", "0110110101101001100110011001100", "0110110101111001100110011001100", 
"0110110110001001100110011001100", "0110110110011001100110011001100", "0110110110101001100110011001100", "0110110110111001100110011001100", 
"0110110111001001100110011001100", "0110110111011001100110011001100", "0110110111101001100110011001100", "0110110111111001100110011001100", 
"0110111000001001100110011001100", "0110111000011001100110011001100", "0110111000101001100110011001100", "0110111000111001100110011001100", 
"0110111001001001100110011001100", "0110111001011001100110011001100", "0110111001101001100110011001100", "0110111001111001100110011001100", 
"0110111010001001100110011001100", "0110111010011001100110011001100", "0110111010101001100110011001100", "0110111010111001100110011001100", 
"0110111011001001100110011001100", "0110111011011001100110011001100", "0110111011101001100110011001100", "0110111011111001100110011001100", 
"0110111100001001100110011001100", "0110111100011001100110011001100", "0110111100101001100110011001100", "0110111100111001100110011001100", 
"0110111101001001100110011001100", "0110111101011001100110011001100", "0110111101101001100110011001100", "0110111101111001100110011001100", 
"0110111110001001100110011001100", "0110111110011001100110011001100", "0110111110101001100110011001100", "0110111110111001100110011001100", 
"0110111111001001100110011001100", "0110111111011001100110011001100", "0110111111101001100110011001100", "0110111111111001100110011001100", 
"0111000000001001100110011001100", "0111000000011001100110011001100", "0111000000101001100110011001100", "0111000000111001100110011001100", 
"0111000001001001100110011001100", "0111000001011001100110011001100", "0111000001101001100110011001100", "0111000001111001100110011001100", 
"0111000010001001100110011001100", "0111000010011001100110011001100", "0111000010101001100110011001100", "0111000010111001100110011001100", 
"0111000011001001100110011001100", "0111000011011001100110011001100", "0111000011101001100110011001100", "0111000011111001100110011001100", 
"0111000100001001100110011001100", "0111000100011001100110011001100", "0111000100101001100110011001100", "0111000100111001100110011001100", 
"0111000101001001100110011001100", "0111000101011001100110011001100", "0111000101101001100110011001100", "0111000101111001100110011001100", 
"0111000110001001100110011001100", "0111000110011001100110011001100", "0111000110101001100110011001100", "0111000110111001100110011001100", 
"0111000111001001100110011001100", "0111000111011001100110011001100", "0111000111101001100110011001100", "0111000111111001100110011001100", 
"0111001000001001100110011001100", "0111001000011001100110011001100", "0111001000101001100110011001100", "0111001000111001100110011001100", 
"0111001001001001100110011001100", "0111001001011001100110011001100", "0111001001101001100110011001100", "0111001001111001100110011001100", 
"0111001010001001100110011001100", "0111001010011001100110011001100", "0111001010101001100110011001100", "0111001010111001100110011001100", 
"0111001011001001100110011001100", "0111001011011001100110011001100", "0111001011101001100110011001100", "0111001011111001100110011001100", 
"0111001100001001100110011001100", "0111001100011001100110011001100", "0111001100101001100110011001100", "0111001100111001100110011001100", 
"0111001101001001100110011001100", "0111001101011001100110011001100", "0111001101101001100110011001100", "0111001101111001100110011001100", 
"0111001110001001100110011001100", "0111001110011001100110011001100", "0111001110101001100110011001100", "0111001110111001100110011001100", 
"0111001111001001100110011001100", "0111001111011001100110011001100", "0111001111101001100110011001100", "0111001111111001100110011001100", 
"0111010000001001100110011001100", "0111010000011001100110011001100", "0111010000101001100110011001100", "0111010000111001100110011001100", 
"0111010001001001100110011001100", "0111010001011001100110011001100", "0111010001101001100110011001100", "0111010001111001100110011001100", 
"0111010010001001100110011001100", "0111010010011001100110011001100", "0111010010101001100110011001100", "0111010010111001100110011001100", 
"0111010011001001100110011001100", "0111010011011001100110011001100", "0111010011101001100110011001100", "0111010011111001100110011001100", 
"0111010100001001100110011001100", "0111010100011001100110011001100", "0111010100101001100110011001100", "0111010100111001100110011001100", 
"0111010101001001100110011001100", "0111010101011001100110011001100", "0111010101101001100110011001100", "0111010101111001100110011001100", 
"0111010110001001100110011001100", "0111010110011001100110011001100", "0111010110101001100110011001100", "0111010110111001100110011001100", 
"0111010111001001100110011001100", "0111010111011001100110011001100", "0111010111101001100110011001100", "0111010111111001100110011001100", 
"0111011000001001100110011001100", "0111011000011001100110011001100", "0111011000101001100110011001100", "0111011000111001100110011001100", 
"0111011001001001100110011001100", "0111011001011001100110011001100", "0111011001101001100110011001100", "0111011001111001100110011001100", 
"0111011010001001100110011001100", "0111011010011001100110011001100", "0111011010101001100110011001100", "0111011010111001100110011001100", 
"0111011011001001100110011001100", "0111011011011001100110011001100", "0111011011101001100110011001100", "0111011011111001100110011001100", 
"0111011100001001100110011001100", "0111011100011001100110011001100", "0111011100101001100110011001100", "0111011100111001100110011001100", 
"0111011101001001100110011001100", "0111011101011001100110011001100", "0111011101101001100110011001100", "0111011101111001100110011001100", 
"0111011110001001100110011001100", "0111011110011001100110011001100", "0111011110101001100110011001100", "0111011110111001100110011001100", 
"0111011111001001100110011001100", "0111011111011001100110011001100", "0111011111101001100110011001100", "0111011111111001100110011001100", 
"0111100000001001100110011001100", "0111100000011001100110011001100", "0111100000101001100110011001100", "0111100000111001100110011001100", 
"0111100001001001100110011001100", "0111100001011001100110011001100", "0111100001101001100110011001100", "0111100001111001100110011001100", 
"0111100010001001100110011001100", "0111100010011001100110011001100", "0111100010101001100110011001100", "0111100010111001100110011001100", 
"0111100011001001100110011001100", "0111100011011001100110011001100", "0111100011101001100110011001100", "0111100011111001100110011001100", 
"0111100100001001100110011001100", "0111100100011001100110011001100", "0111100100101001100110011001100", "0111100100111001100110011001100", 
"0111100101001001100110011001100", "0111100101011001100110011001100", "0111100101101001100110011001100", "0111100101111001100110011001100", 
"0111100110001001100110011001100", "0111100110011001100110011001100", "0111100110101001100110011001100", "0111100110111001100110011001100", 
"0111100111001001100110011001100", "0111100111011001100110011001100", "0111100111101001100110011001100", "0111100111111001100110011001100", 
"0111101000001001100110011001100", "0111101000011001100110011001100", "0111101000101001100110011001100", "0111101000111001100110011001100", 
"0111101001001001100110011001100", "0111101001011001100110011001100", "0111101001101001100110011001100", "0111101001111001100110011001100", 
"0111101010001001100110011001100", "0111101010011001100110011001100", "0111101010101001100110011001100", "0111101010111001100110011001100", 
"0111101011001001100110011001100", "0111101011011001100110011001100", "0111101011101001100110011001100", "0111101011111001100110011001100", 
"0111101100001001100110011001100", "0111101100011001100110011001100", "0111101100101001100110011001100", "0111101100111001100110011001100", 
"0111101101001001100110011001100", "0111101101011001100110011001100", "0111101101101001100110011001100", "0111101101111001100110011001100", 
"0111101110001001100110011001100", "0111101110011001100110011001100", "0111101110101001100110011001100", "0111101110111001100110011001100", 
"0111101111001001100110011001100", "0111101111011001100110011001100", "0111101111101001100110011001100", "0111101111111001100110011001100", 
"0111110000001001100110011001100", "0111110000011001100110011001100", "0111110000101001100110011001100", "0111110000111001100110011001100", 
"0111110001001001100110011001100", "0111110001011001100110011001100", "0111110001101001100110011001100", "0111110001111001100110011001100", 
"0111110010001001100110011001100", "0111110010011001100110011001100", "0111110010101001100110011001100", "0111110010111001100110011001100", 
"0111110011001001100110011001100", "0111110011011001100110011001100", "0111110011101001100110011001100", "0111110011111001100110011001100", 
"0111110100001001100110011001100", "0111110100011001100110011001100", "0111110100101001100110011001100", "0111110100111001100110011001100", 
"0111110101001001100110011001100", "0111110101011001100110011001100", "0111110101101001100110011001100", "0111110101111001100110011001100", 
"0111110110001001100110011001100", "0111110110011001100110011001100", "0111110110101001100110011001100", "0111110110111001100110011001100", 
"0111110111001001100110011001100", "0111110111011001100110011001100", "0111110111101001100110011001100", "0111110111111001100110011001100", 
"0111111000001001100110011001100", "0111111000011001100110011001100", "0111111000101001100110011001100", "0111111000111001100110011001100", 
"0111111001001001100110011001100", "0111111001011001100110011001100", "0111111001101001100110011001100", "0111111001111001100110011001100", 
"0111111010001001100110011001100", "0111111010011001100110011001100", "0111111010101001100110011001100", "0111111010111001100110011001100", 
"0111111011001001100110011001100", "0111111011011001100110011001100", "0111111011101001100110011001100", "0111111011111001100110011001100", 
"0111111100001001100110011001100", "0111111100011001100110011001100", "0111111100101001100110011001100", "0111111100111001100110011001100", 
"0111111101001001100110011001100", "0111111101011001100110011001100", "0111111101101001100110011001100", "0111111101111001100110011001100", 
"0111111110001001100110011001100", "0111111110011001100110011001100", "0111111110101001100110011001100", "0111111110111001100110011001100", 
"0111111111001001100110011001100", "0111111111011001100110011001100", "0111111111101001100110011001100", "0111111111111001100110011001100"
);
type muon_pt_lut_sfixed_array is array (0 to 2**(D_S_I_MUON_V2.pt_high-D_S_I_MUON_V2.pt_low+1)-1) of sfixed(8 downto -20);
constant MU_PT_LUT_SFIXED : muon_pt_lut_sfixed_array := (
"00000000000000000000000000000", "00000000001001100110011001100", "00000000011001100110011001100", "00000000101001100110011001100", 
"00000000111001100110011001100", "00000001001001100110011001100", "00000001011001100110011001100", "00000001101001100110011001100", 
"00000001111001100110011001100", "00000010001001100110011001100", "00000010011001100110011001100", "00000010101001100110011001100", 
"00000010111001100110011001100", "00000011001001100110011001100", "00000011011001100110011001100", "00000011101001100110011001100", 
"00000011111001100110011001100", "00000100001001100110011001100", "00000100011001100110011001100", "00000100101001100110011001100", 
"00000100111001100110011001100", "00000101001001100110011001100", "00000101011001100110011001100", "00000101101001100110011001100", 
"00000101111001100110011001100", "00000110001001100110011001100", "00000110011001100110011001100", "00000110101001100110011001100", 
"00000110111001100110011001100", "00000111001001100110011001100", "00000111011001100110011001100", "00000111101001100110011001100", 
"00000111111001100110011001100", "00001000001001100110011001100", "00001000011001100110011001100", "00001000101001100110011001100", 
"00001000111001100110011001100", "00001001001001100110011001100", "00001001011001100110011001100", "00001001101001100110011001100", 
"00001001111001100110011001100", "00001010001001100110011001100", "00001010011001100110011001100", "00001010101001100110011001100", 
"00001010111001100110011001100", "00001011001001100110011001100", "00001011011001100110011001100", "00001011101001100110011001100", 
"00001011111001100110011001100", "00001100001001100110011001100", "00001100011001100110011001100", "00001100101001100110011001100", 
"00001100111001100110011001100", "00001101001001100110011001100", "00001101011001100110011001100", "00001101101001100110011001100", 
"00001101111001100110011001100", "00001110001001100110011001100", "00001110011001100110011001100", "00001110101001100110011001100", 
"00001110111001100110011001100", "00001111001001100110011001100", "00001111011001100110011001100", "00001111101001100110011001100", 
"00001111111001100110011001100", "00010000001001100110011001100", "00010000011001100110011001100", "00010000101001100110011001100", 
"00010000111001100110011001100", "00010001001001100110011001100", "00010001011001100110011001100", "00010001101001100110011001100", 
"00010001111001100110011001100", "00010010001001100110011001100", "00010010011001100110011001100", "00010010101001100110011001100", 
"00010010111001100110011001100", "00010011001001100110011001100", "00010011011001100110011001100", "00010011101001100110011001100", 
"00010011111001100110011001100", "00010100001001100110011001100", "00010100011001100110011001100", "00010100101001100110011001100", 
"00010100111001100110011001100", "00010101001001100110011001100", "00010101011001100110011001100", "00010101101001100110011001100", 
"00010101111001100110011001100", "00010110001001100110011001100", "00010110011001100110011001100", "00010110101001100110011001100", 
"00010110111001100110011001100", "00010111001001100110011001100", "00010111011001100110011001100", "00010111101001100110011001100", 
"00010111111001100110011001100", "00011000001001100110011001100", "00011000011001100110011001100", "00011000101001100110011001100", 
"00011000111001100110011001100", "00011001001001100110011001100", "00011001011001100110011001100", "00011001101001100110011001100", 
"00011001111001100110011001100", "00011010001001100110011001100", "00011010011001100110011001100", "00011010101001100110011001100", 
"00011010111001100110011001100", "00011011001001100110011001100", "00011011011001100110011001100", "00011011101001100110011001100", 
"00011011111001100110011001100", "00011100001001100110011001100", "00011100011001100110011001100", "00011100101001100110011001100", 
"00011100111001100110011001100", "00011101001001100110011001100", "00011101011001100110011001100", "00011101101001100110011001100", 
"00011101111001100110011001100", "00011110001001100110011001100", "00011110011001100110011001100", "00011110101001100110011001100", 
"00011110111001100110011001100", "00011111001001100110011001100", "00011111011001100110011001100", "00011111101001100110011001100", 
"00011111111001100110011001100", "00100000001001100110011001100", "00100000011001100110011001100", "00100000101001100110011001100", 
"00100000111001100110011001100", "00100001001001100110011001100", "00100001011001100110011001100", "00100001101001100110011001100", 
"00100001111001100110011001100", "00100010001001100110011001100", "00100010011001100110011001100", "00100010101001100110011001100", 
"00100010111001100110011001100", "00100011001001100110011001100", "00100011011001100110011001100", "00100011101001100110011001100", 
"00100011111001100110011001100", "00100100001001100110011001100", "00100100011001100110011001100", "00100100101001100110011001100", 
"00100100111001100110011001100", "00100101001001100110011001100", "00100101011001100110011001100", "00100101101001100110011001100", 
"00100101111001100110011001100", "00100110001001100110011001100", "00100110011001100110011001100", "00100110101001100110011001100", 
"00100110111001100110011001100", "00100111001001100110011001100", "00100111011001100110011001100", "00100111101001100110011001100", 
"00100111111001100110011001100", "00101000001001100110011001100", "00101000011001100110011001100", "00101000101001100110011001100", 
"00101000111001100110011001100", "00101001001001100110011001100", "00101001011001100110011001100", "00101001101001100110011001100", 
"00101001111001100110011001100", "00101010001001100110011001100", "00101010011001100110011001100", "00101010101001100110011001100", 
"00101010111001100110011001100", "00101011001001100110011001100", "00101011011001100110011001100", "00101011101001100110011001100", 
"00101011111001100110011001100", "00101100001001100110011001100", "00101100011001100110011001100", "00101100101001100110011001100", 
"00101100111001100110011001100", "00101101001001100110011001100", "00101101011001100110011001100", "00101101101001100110011001100", 
"00101101111001100110011001100", "00101110001001100110011001100", "00101110011001100110011001100", "00101110101001100110011001100", 
"00101110111001100110011001100", "00101111001001100110011001100", "00101111011001100110011001100", "00101111101001100110011001100", 
"00101111111001100110011001100", "00110000001001100110011001100", "00110000011001100110011001100", "00110000101001100110011001100", 
"00110000111001100110011001100", "00110001001001100110011001100", "00110001011001100110011001100", "00110001101001100110011001100", 
"00110001111001100110011001100", "00110010001001100110011001100", "00110010011001100110011001100", "00110010101001100110011001100", 
"00110010111001100110011001100", "00110011001001100110011001100", "00110011011001100110011001100", "00110011101001100110011001100", 
"00110011111001100110011001100", "00110100001001100110011001100", "00110100011001100110011001100", "00110100101001100110011001100", 
"00110100111001100110011001100", "00110101001001100110011001100", "00110101011001100110011001100", "00110101101001100110011001100", 
"00110101111001100110011001100", "00110110001001100110011001100", "00110110011001100110011001100", "00110110101001100110011001100", 
"00110110111001100110011001100", "00110111001001100110011001100", "00110111011001100110011001100", "00110111101001100110011001100", 
"00110111111001100110011001100", "00111000001001100110011001100", "00111000011001100110011001100", "00111000101001100110011001100", 
"00111000111001100110011001100", "00111001001001100110011001100", "00111001011001100110011001100", "00111001101001100110011001100", 
"00111001111001100110011001100", "00111010001001100110011001100", "00111010011001100110011001100", "00111010101001100110011001100", 
"00111010111001100110011001100", "00111011001001100110011001100", "00111011011001100110011001100", "00111011101001100110011001100", 
"00111011111001100110011001100", "00111100001001100110011001100", "00111100011001100110011001100", "00111100101001100110011001100", 
"00111100111001100110011001100", "00111101001001100110011001100", "00111101011001100110011001100", "00111101101001100110011001100", 
"00111101111001100110011001100", "00111110001001100110011001100", "00111110011001100110011001100", "00111110101001100110011001100", 
"00111110111001100110011001100", "00111111001001100110011001100", "00111111011001100110011001100", "00111111101001100110011001100", 
"00111111111001100110011001100", "01000000001001100110011001100", "01000000011001100110011001100", "01000000101001100110011001100", 
"01000000111001100110011001100", "01000001001001100110011001100", "01000001011001100110011001100", "01000001101001100110011001100", 
"01000001111001100110011001100", "01000010001001100110011001100", "01000010011001100110011001100", "01000010101001100110011001100", 
"01000010111001100110011001100", "01000011001001100110011001100", "01000011011001100110011001100", "01000011101001100110011001100", 
"01000011111001100110011001100", "01000100001001100110011001100", "01000100011001100110011001100", "01000100101001100110011001100", 
"01000100111001100110011001100", "01000101001001100110011001100", "01000101011001100110011001100", "01000101101001100110011001100", 
"01000101111001100110011001100", "01000110001001100110011001100", "01000110011001100110011001100", "01000110101001100110011001100", 
"01000110111001100110011001100", "01000111001001100110011001100", "01000111011001100110011001100", "01000111101001100110011001100", 
"01000111111001100110011001100", "01001000001001100110011001100", "01001000011001100110011001100", "01001000101001100110011001100", 
"01001000111001100110011001100", "01001001001001100110011001100", "01001001011001100110011001100", "01001001101001100110011001100", 
"01001001111001100110011001100", "01001010001001100110011001100", "01001010011001100110011001100", "01001010101001100110011001100", 
"01001010111001100110011001100", "01001011001001100110011001100", "01001011011001100110011001100", "01001011101001100110011001100", 
"01001011111001100110011001100", "01001100001001100110011001100", "01001100011001100110011001100", "01001100101001100110011001100", 
"01001100111001100110011001100", "01001101001001100110011001100", "01001101011001100110011001100", "01001101101001100110011001100", 
"01001101111001100110011001100", "01001110001001100110011001100", "01001110011001100110011001100", "01001110101001100110011001100", 
"01001110111001100110011001100", "01001111001001100110011001100", "01001111011001100110011001100", "01001111101001100110011001100", 
"01001111111001100110011001100", "01010000001001100110011001100", "01010000011001100110011001100", "01010000101001100110011001100", 
"01010000111001100110011001100", "01010001001001100110011001100", "01010001011001100110011001100", "01010001101001100110011001100", 
"01010001111001100110011001100", "01010010001001100110011001100", "01010010011001100110011001100", "01010010101001100110011001100", 
"01010010111001100110011001100", "01010011001001100110011001100", "01010011011001100110011001100", "01010011101001100110011001100", 
"01010011111001100110011001100", "01010100001001100110011001100", "01010100011001100110011001100", "01010100101001100110011001100", 
"01010100111001100110011001100", "01010101001001100110011001100", "01010101011001100110011001100", "01010101101001100110011001100", 
"01010101111001100110011001100", "01010110001001100110011001100", "01010110011001100110011001100", "01010110101001100110011001100", 
"01010110111001100110011001100", "01010111001001100110011001100", "01010111011001100110011001100", "01010111101001100110011001100", 
"01010111111001100110011001100", "01011000001001100110011001100", "01011000011001100110011001100", "01011000101001100110011001100", 
"01011000111001100110011001100", "01011001001001100110011001100", "01011001011001100110011001100", "01011001101001100110011001100", 
"01011001111001100110011001100", "01011010001001100110011001100", "01011010011001100110011001100", "01011010101001100110011001100", 
"01011010111001100110011001100", "01011011001001100110011001100", "01011011011001100110011001100", "01011011101001100110011001100", 
"01011011111001100110011001100", "01011100001001100110011001100", "01011100011001100110011001100", "01011100101001100110011001100", 
"01011100111001100110011001100", "01011101001001100110011001100", "01011101011001100110011001100", "01011101101001100110011001100", 
"01011101111001100110011001100", "01011110001001100110011001100", "01011110011001100110011001100", "01011110101001100110011001100", 
"01011110111001100110011001100", "01011111001001100110011001100", "01011111011001100110011001100", "01011111101001100110011001100", 
"01011111111001100110011001100", "01100000001001100110011001100", "01100000011001100110011001100", "01100000101001100110011001100", 
"01100000111001100110011001100", "01100001001001100110011001100", "01100001011001100110011001100", "01100001101001100110011001100", 
"01100001111001100110011001100", "01100010001001100110011001100", "01100010011001100110011001100", "01100010101001100110011001100", 
"01100010111001100110011001100", "01100011001001100110011001100", "01100011011001100110011001100", "01100011101001100110011001100", 
"01100011111001100110011001100", "01100100001001100110011001100", "01100100011001100110011001100", "01100100101001100110011001100", 
"01100100111001100110011001100", "01100101001001100110011001100", "01100101011001100110011001100", "01100101101001100110011001100", 
"01100101111001100110011001100", "01100110001001100110011001100", "01100110011001100110011001100", "01100110101001100110011001100", 
"01100110111001100110011001100", "01100111001001100110011001100", "01100111011001100110011001100", "01100111101001100110011001100", 
"01100111111001100110011001100", "01101000001001100110011001100", "01101000011001100110011001100", "01101000101001100110011001100", 
"01101000111001100110011001100", "01101001001001100110011001100", "01101001011001100110011001100", "01101001101001100110011001100", 
"01101001111001100110011001100", "01101010001001100110011001100", "01101010011001100110011001100", "01101010101001100110011001100", 
"01101010111001100110011001100", "01101011001001100110011001100", "01101011011001100110011001100", "01101011101001100110011001100", 
"01101011111001100110011001100", "01101100001001100110011001100", "01101100011001100110011001100", "01101100101001100110011001100", 
"01101100111001100110011001100", "01101101001001100110011001100", "01101101011001100110011001100", "01101101101001100110011001100", 
"01101101111001100110011001100", "01101110001001100110011001100", "01101110011001100110011001100", "01101110101001100110011001100", 
"01101110111001100110011001100", "01101111001001100110011001100", "01101111011001100110011001100", "01101111101001100110011001100", 
"01101111111001100110011001100", "01110000001001100110011001100", "01110000011001100110011001100", "01110000101001100110011001100", 
"01110000111001100110011001100", "01110001001001100110011001100", "01110001011001100110011001100", "01110001101001100110011001100", 
"01110001111001100110011001100", "01110010001001100110011001100", "01110010011001100110011001100", "01110010101001100110011001100", 
"01110010111001100110011001100", "01110011001001100110011001100", "01110011011001100110011001100", "01110011101001100110011001100", 
"01110011111001100110011001100", "01110100001001100110011001100", "01110100011001100110011001100", "01110100101001100110011001100", 
"01110100111001100110011001100", "01110101001001100110011001100", "01110101011001100110011001100", "01110101101001100110011001100", 
"01110101111001100110011001100", "01110110001001100110011001100", "01110110011001100110011001100", "01110110101001100110011001100", 
"01110110111001100110011001100", "01110111001001100110011001100", "01110111011001100110011001100", "01110111101001100110011001100", 
"01110111111001100110011001100", "01111000001001100110011001100", "01111000011001100110011001100", "01111000101001100110011001100", 
"01111000111001100110011001100", "01111001001001100110011001100", "01111001011001100110011001100", "01111001101001100110011001100", 
"01111001111001100110011001100", "01111010001001100110011001100", "01111010011001100110011001100", "01111010101001100110011001100", 
"01111010111001100110011001100", "01111011001001100110011001100", "01111011011001100110011001100", "01111011101001100110011001100", 
"01111011111001100110011001100", "01111100001001100110011001100", "01111100011001100110011001100", "01111100101001100110011001100", 
"01111100111001100110011001100", "01111101001001100110011001100", "01111101011001100110011001100", "01111101101001100110011001100", 
"01111101111001100110011001100", "01111110001001100110011001100", "01111110011001100110011001100", "01111110101001100110011001100", 
"01111110111001100110011001100", "01111111001001100110011001100", "01111111011001100110011001100", "01111111101001100110011001100"
);
type calo_calo_diff_eta_lut_sfixed_array is array (0 to 2**MAX_CALO_ETA_BITS-1) of sfixed(4 downto -20);
constant CALO_CALO_DIFF_ETA_LUT_SFIXED : calo_calo_diff_eta_lut_sfixed_array := (
"0000000000000000000000000", "0000000001011010000111000", "0000000010110010001011010", "0000000100001100010010010", 
"0000000101100100010110100", "0000000110111100011010100", "0000001000010110100001110", "0000001001110000101000110", 
"0000001011001000101101000", "0000001100100000110001000", "0000001101111010111000010", "0000001111010100111111010", 
"0000010000101101000011100", "0000010010000111001010110", "0000010011011111001110110", "0000010100111001010110000", 
"0000010110010001011010000", "0000010111101001011110000", "0000011001000011100101010", "0000011010011011101001010", 
"0000011011110101110000100", "0000011101001111110111110", "0000011110100111111011110", "0000100000000010000011000", 
"0000100001011010000111000", "0000100010110100001110010", "0000100100001100010010010", "0000100101100100010110100", 
"0000100110111110011101100", "0000101000010110100001110", "0000101001110000101000110", "0000101011001000101101000", 
"0000101100100010110100000", "0000101101111100111011010", "0000101111010100111111010", "0000110000101111000110100", 
"0000110010000111001010110", "0000110011100001010001110", "0000110100111001010110000", "0000110110010011011101000", 
"0000110111101011100001010", "0000111001000011100101010", "0000111010011101101100100", "0000111011110101110000100", 
"0000111101001111110111110", "0000111110100111111011110", "0001000000000010000011000", "0001000001011010000111000", 
"0001000010110100001110010", "0001000100001110010101100", "0001000101100110011001100", "0001000110111110011101100", 
"0001001000011000100100110", "0001001001110010101100000", "0001001011001010110000000", "0001001100100010110100000", 
"0001001101111100111011010", "0001001111010111000010100", "0001010000101111000110100", "0001010010001001001101110", 
"0001010011100001010001110", "0001010100111001010110000", "0001010110010011011101000", "0001010111101101100100010", 
"0001011001000101101000010", "0001011010011101101100100", "0001011011110111110011100", "0001011101010001111010110", 
"0001011110101001111110110", "0001100000000010000011000", "0001100001011100001010000", "0001100010110110010001010", 
"0001100100001110010101100", "0001100101101000011100100", "0001100111000000100000110", "0001101000011000100100110", 
"0001101001110010101100000", "0001101011001100110011000", "0001101100100100110111010", "0001101101111100111011010", 
"0001101111010111000010100", "0001110000110001001001100", "0001110010001001001101110", "0001110011100001010001110", 
"0001110100111011011001000", "0001110110010101100000010", "0001110111101101100100010", "0001111001000101101000010", 
"0001111010011111101111100", "0001111011110111110011100", "0001111101010001111010110", "0001111110101100000010000", 
"0010000000000100000110000", "0010000001011100001010000", "0010000010110110010001010", "0010000100001110010101100", 
"0010000101101000011100100", "0010000111000010100011110", "0010001000011010100111110", "0010001001110100101111000", 
"0010001011001100110011000", "0010001100100100110111010", "0010001101111110111110010", "0010001111010111000010100", 
"0010010000110001001001100", "0010010010001011010000110", "0010010011100011010100110", "0010010100111101011100000", 
"0010010110010101100000010", "0010010111101101100100010", "0010011001000111101011100", "0010011010100001110010100", 
"0010011011111001110110110", "0010011101010011111101110", "0010011110101100000010000", "0010100000000100000110000", 
"0010100001011110001101010", "0010100010110110010001010", "0010100100010000011000100", "0010100101101010011111100", 
"0010100111000010100011110", "0010101000011100101011000", "0010101001110100101111000", "0010101011001100110011000", 
"0010101100100110111010010", "0010101110000001000001100", "0010101111011001000101100", "0010110000110011001100110", 
"0010110010001011010000110", "0010110011100011010100110", "0010110100111101011100000", "0010110110010101100000010", 
"0010110111101111100111010", "0010111001001001101110100", "0010111010100001110010100", "0010111011111011111001110", 
"0010111101010011111101110", "0010111110101100000010000", "0011000000000110001001000", "0011000001100000010000010", 
"0011000010111000010100010", "0011000100010010011011100", "0011000101101010011111100", "0011000111000010100011110", 
"0011001000011100101011000", "0011001001110100101111000", "0011001011001110110110010", "0011001100101000111101010", 
"0011001110000001000001100", "0011001111011011001000100", "0011010000110011001100110", "0011010010001011010000110", 
"0011010011100101011000000", "0011010100111111011111000", "0011010110010111100011010", "0011010111110001101010010", 
"0011011001001001101110100", "0011011010100001110010100", "0011011011111011111001110", "0011011101010011111101110", 
"0011011110101110000101000", "0011100000001000001100010", "0011100001100000010000010", "0011100010111010010111100", 
"0011100100010010011011100", "0011100101101010011111100", "0011100111000100100110110", "0011101000011100101011000", 
"0011101001110110110010000", "0011101011010000111001010", "0011101100101000111101010", "0011101110000001000001100", 
"0011101111011011001000100", "0011110000110011001100110", "0011110010001101010011110", "0011110011100111011011000", 
"0011110100111111011111000", "0011110110011001100110010", "0011110111110001101010010", "0011111001001001101110100", 
"0011111010100011110101110", "0011111011111011111001110", "0011111101010110000001000", "0011111110110000001000000", 
"0100000000001000001100010", "0100000001100000010000010", "0100000010111010010111100", "0100000100010010011011100", 
"0100000101101100100010110", "0100000111000100100110110", "0100001000011110101110000", "0100001001110110110010000", 
"0100001011010000111001010", "0100001100101011000000100", "0100001110000011000100100", "0100001111011101001011110", 
"0100010000110101001111110", "0100010010001111010111000", "0100010011100111011011000", "0100010101000001100010010", 
"0100010110011001100110010", "0100010111110011101101100", "0100011001001011110001100", "0100011010100011110101110", 
"0100011011111101111100110", "0100011101010110000001000", "0100011110110000001000000", "0100100000001010001111010", 
"0100100001100010010011010", "0100100010111100011010100", "0100100100010100011110100", "0100100101101110100101110", 
"0100100111000110101001110", "0100101000100000110001000", "0100101001111000110101000", "0100101011010010111100010", 
"0100101100101011000000100", "0100101110000011000100100", "0100101111011101001011110", "0100110000110101001111110", 
"0100110010001111010111000", "0100110011101001011110000", "0100110101000001100010010", "0100110110011011101001010", 
"0100110111110011101101100", "0100111001001101110100100", "0100111010100101111000110", "0100111011111111111111110", 
"0100111101011000000100000", "0100111110110010001011010", "0000000000000000000000000", "0000000000000000000000000", 
"0000000000000000000000000", "0000000000000000000000000", "0000000000000000000000000", "0000000000000000000000000", 
"0000000000000000000000000", "0000000000000000000000000", "0000000000000000000000000", "0000000000000000000000000", 
"0000000000000000000000000", "0000000000000000000000000", "0000000000000000000000000", "0000000000000000000000000", 
"0000000000000000000000000", "0000000000000000000000000", "0000000000000000000000000", "0000000000000000000000000", 
"0000000000000000000000000", "0000000000000000000000000", "0000000000000000000000000", "0000000000000000000000000", 
"0000000000000000000000000", "0000000000000000000000000", "0000000000000000000000000", "0000000000000000000000000"
);
type calo_calo_diff_phi_lut_sfixed_array is array (0 to 2**MAX_CALO_PHI_BITS-1) of sfixed(3 downto -20);
constant CALO_CALO_DIFF_PHI_LUT_SFIXED : calo_calo_diff_phi_lut_sfixed_array := (
"000000000000000000000000", "000000001011010000111000", "000000010110010001011010", "000000100001100010010010", 
"000000101100110011001100", "000000110111110011101100", "000001000011000100100110", "000001001110000101000110", 
"000001011001010110000000", "000001100100100110111010", "000001101111100111011010", "000001111010111000010100", 
"000010000110001001001100", "000010010001001001101110", "000010011100011010100110", "000010100111011011001000", 
"000010110010101100000010", "000010111101111100111010", "000011001000111101011100", "000011010100001110010100", 
"000011011111011111001110", "000011101010011111101110", "000011110101110000101000", "000100000001000001100010", 
"000100001100000010000010", "000100010111010010111100", "000100100010010011011100", "000100101101100100010110", 
"000100111000110101001110", "000101000011110101110000", "000101001111000110101000", "000101011010010111100010", 
"000101100101011000000100", "000101110000101000111100", "000101111011111001110110", "000110000110111010010110", 
"000110010010001011010000", "000110011101001011110000", "000110101000011100101010", "000110110011101101100100", 
"000110111110101110000100", "000111001001111110111110", "000111010101001111110110", "000111100000010000011000", 
"000111101011100001010000", "000111110110100001110010", "001000000001110010101100", "001000001101000011100100", 
"001000011000000100000110", "001000100011010100111110", "001000101110100101111000", "001000111001100110011000", 
"001001000100110111010010", "001001010000001000001100", "001001011011001000101100", "001001100110011001100110", 
"001001110001011010000110", "001001111100101011000000", "001010000111111011111000", "001010010010111100011010", 
"001010011110001101010010", "001010101001011110001100", "001010110100011110101110", "001010111111101111100110", 
"001011001011000000100000", "001011010110000001000000", "001011100001010001111010", "001011101100010010011010", 
"001011110111100011010100", "001100000010110100001110", "001100001101110100101110", "001100011001000101101000", 
"001100100100010110100000", "001100101111010111000010", "001100111010100111111010", "001101000101101000011100", 
"001101010000111001010110", "001101011100001010001110", "001101100111001010110000", "001101110010011011101000", 
"001101111101101100100010", "001110001000101101000010", "001110010011111101111100", "001110011111001110110110", 
"001110101010001111010110", "001110110101100000010000", "001111000000100000110000", "001111001011110001101010", 
"001111010111000010100010", "001111100010000011000100", "001111101101010011111100", "001111111000100100110110", 
"010000000011100101011000", "010000001110110110010000", "010000011010000111001010", "010000100101000111101010", 
"010000110000011000100100", "010000111011011001000100", "010001000110101001111110", "010001010001111010111000", 
"010001011100111011011000", "010001101000001100010010", "010001110011011101001010", "010001111110011101101100", 
"010010001001101110100100", "010010010100101111000110", "010010011111111111111110", "010010101011010000111000", 
"010010110110010001011010", "010011000001100010010010", "010011001100110011001100", "010011010111110011101100", 
"010011100011000100100110", "010011101110010101100000", "010011111001010110000000", "010100000100100110111010", 
"010100001111100111011010", "010100011010111000010100", "010100100110001001001100", "010100110001001001101110", 
"010100111100011010100110", "010101000111101011100000", "010101010010101100000010", "010101011101111100111010", 
"010101101001001101110100", "010101110100001110010100", "010101111111011111001110", "010110001010011111101110", 
"010110010101110000101000", "010110100001000001100010", "010110101100000010000010", "010110110111010010111100", 
"010111000010100011110100", "010111001101100100010110", "010111011000110101001110", "010111100011110101110000", 
"010111101111000110101000", "010111111010010111100010", "011000000101011000000100", "011000010000101000111100", 
"011000011011111001110110", "011000100110111010010110", "011000110010001011010000", "011000111101011100001010", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000"
);
type calo_calo_cosh_deta_lut_sfixed_array is array (0 to 2**MAX_CALO_ETA_BITS-1) of sfixed(14 downto -20);
constant CALO_CALO_COSH_DETA_LUT_SFIXED : calo_calo_cosh_deta_lut_sfixed_array := (
"00000000000000100000000000000000000", "00000000000000100000000010000011000", "00000000000000100000001000001100010", "00000000000000100000010010011011100", 
"00000000000000100000011110101110000", "00000000000000100000110001001001100", "00000000000000100001000101101000010", "00000000000000100001100000010000010", 
"00000000000000100001111100111011010", "00000000000000100010011111101111100", "00000000000000100011000100100110110", "00000000000000100011101111100111010", 
"00000000000000100100011100101011000", "00000000000000100101001111110111110", "00000000000000100110000111001010110", "00000000000000100111000100100110110", 
"00000000000000101000000100000110000", "00000000000000101001001001101110100", "00000000000000101010010101100000010", "00000000000000101011100011010100110", 
"00000000000000101100111001010110000", "00000000000000101110010011011101000", "00000000000000101111110011101101100", "00000000000000110001011010000111000", 
"00000000000000110011000100100110110", "00000000000000110100110111010010110", "00000000000000110110110000001000000", "00000000000000111000101111000110100", 
"00000000000000111010110100001110010", "00000000000000111101000001100010010", "00000000000000111111010100111111010", "00000000000001000001110010101100000", 
"00000000000001000100010110100001110", "00000000000001000111000010100011110", "00000000000001001001110110110010000", "00000000000001001100110101001111110", 
"00000000000001001111111011111001110", "00000000000001010011001100110011000", "00000000000001010110100111111011110", "00000000000001011010001101010011110", 
"00000000000001011101111100111011010", "00000000000001100001111000110101000", "00000000000001100110000001000001100", "00000000000001101010010101100000010", 
"00000000000001101110110110010001010", "00000000000001110011100011010100110", "00000000000001111000100000110001000", "00000000000001111101101010011111100", 
"00000000000010000011000100100110110", "00000000000010001000101111000110100", "00000000000010001110101001111110110", "00000000000010010100110101001111110", 
"00000000000010011011010010111100010", "00000000000010100010000011000100100", "00000000000010101001000111101011100", "00000000000010110000100000110001000", 
"00000000000010111000001110010101100", "00000000000011000000010100011110100", "00000000000011001000101111000110100", "00000000000011010001100010010011010", 
"00000000000011011010110000001000000", "00000000000011100100011000100100110", "00000000000011101110011011101001010", "00000000000011111000111101011100000", 
"00000000000100000011111011111001110", "00000000000100001111011001000101100", "00000000000100011011011001000101100", "00000000000100100111111001110110110", 
"00000000000100110100111111011111000", "00000000000101000010101001111110110", "00000000000101010000111011011001000", "00000000000101011111110101110000100", 
"00000000000101101111011011001000100", "00000000000101111111101011100001010", "00000000000110010000101101000011100", "00000000000110100010011101101100100", 
"00000000000110110100111111011111000", "00000000000111001000011000100100110", "00000000000111011100100110111010010", "00000000000111110001110000101000110", 
"00000000001000000111110101110000100", "00000000001000011110111010010111100", "00000000001000110111000000100000110", "00000000001001010000001100010010010", 
"00000000001001101010011101101100100", "00000000001010000101111100111011010", "00000000001010100010100111111011110", "00000000001011000000100100110111010", 
"00000000001011011111110111110011100", "00000000001100000000100100110111010", "00000000001100100010101110000101000", "00000000001101000110010111100011010", 
"00000000001101101011100111011011000", "00000000001110010010100001110010100", "00000000001110111011001000101101000", "00000000001111100101100110011001100", 
"00000000010000010001111010111000010", "00000000010001000000001110010101100", "00000000010001110000100100110111010", "00000000010010100011000110101001110", 
"00000000010011010111110111110011100", "00000000010100001110111110011101100", "00000000010101001000100000110001000", "00000000010110000100101000111101010", 
"00000000010111000011011011001000100", "00000000011000000101000001100010010", "00000000011001001001100000010000010", "00000000011010010001000011100101010", 
"00000000011011011011110001101010010", "00000000011100101001110100101111000", "00000000011101111011010111000010100", "00000000011111010000100000110001000", 
"00000000100000101001011100001010000", "00000000100010000110010011011101000", "00000000100011100111010100111111010", "00000000100101001100101011000000100", 
"00000000100110110110011111101111100", "00000000101000100101000001100010010", "00000000101010011000011110101110000", "00000000101100010001000101101000010", 
"00000000101110001111000010100011110", "00000000110000010010100101111000110", "00000000110010011011111111111111110", "00000000110100101011011111001110110", 
"00000000110111000001011000000100000", "00000000111001011101111100111011010", "00000000111100000001011100001010000", "00000000111110101100001110010101100", 
"00000001000001011110100111111011110", "00000001000100011000111011011001000", "00000001000111011011100001010001110", "00000001001010100110110000001000000", 
"00000001001101111011000010100011110", "00000001010001011000110001001001100", "00000001010101000000010110100001110", "00000001011000110010001101010011110", 
"00000001011100101110110110010001010", "00000001100000110110101100000010000", "00000001100101001010010011011101000", "00000001101001101010001001001101110", 
"00000001101110010110110010001011010", "00000001110011010000110011001100110", "00000001111000011000110001001001100", "00000001111101101111010010111100010", 
"00000010000011010101000101101000010", "00000010001001001010110010001011010", "00000010001111010001000101101000010", "00000010010101101000101111000110100", 
"00000010011100010010011111101111100", "00000010100011001111001110110110010", "00000010101010011111101101100100010", "00000010110010000100110101001111110", 
"00000010111001111111100001010001110", "00000011000010010000110001001001100", "00000011001010111001100010010011010", "00000011010011111010110110010001010", 
"00000011011101010101110110110010000", "00000011100111001011101011100001010", "00000011110001011101011110001101010", "00000011111100001100100010110100000", 
"00000100000111011010001001001101110", "00000100010011000111101011100001010", "00000100011111010110011111101111100", "00000100101100001000001000001100010", 
"00000100111001011110001001001101110", "00000101000111011010000101000111100", "00000101010101111101101100100010110", "00000101100101001010110000001000000", 
"00000101110101000011000010100011110", "00000110000101101000100010110100000", "00000110010110111101001101110100100", "00000110101001000011001010110000000", 
"00000110111011111100101000111101010", "00000111001111101011110101110000100", "00000111100100010011001110110110010", "00000111111001110101010001111010110", 
"00001000010000010100100110111010010", "00001000100111110011111001110110110", "00001001000000010110000011000100100", "00001001011001111110000001000001100", 
"00001001110100101110111000010100010", "00001010010000101011111001110110110", "00001010101101111000011100101011000", "00001011001100011000000110001001000", 
"00001011101100001110011111101111100", "00001100001101011111100001010001110", "00001100110000001111001110110110010", "00001101010100100001110000101000110", 
"00001101111010011011100101011000000", "00001110100010000001001111110111110", "00001111001011010111100101011000000", "00001111110110100011100011010100110", 
"00010000100011101010011001100110010", "00010001010010110001100110011001100", "00010010000011111110110110010001010", "00010010110111011000001000001100010", 
"00010011101101000011101001011110000", "00010100100101000111111011111001110", "00010101011111101011101101100100010", "00010110011100110110001001001101110", 
"00010111011100101110100101111000110", "00011000011111011100110101001111110", "00011001100101001000111011011001000", "00011010101101111011010010111100010", 
"00011011111001111100110011001100110", "00011101001001010110100101111000110", "00011110011100010010010101100000010", "00011111110010111010000101000111100", 
"00100001001101011000010010011011100", "00100010101011110111111011111001110", "00100100001110100100011100101011000", "00100101110101101001110010101100000", 
"00100111100001010100011100101011000", "00101001010001110001011110001101010", "00101011000111001110011111101111100", "00101101000001111001101100100010110", 
"00101111000010000001111110111110010", "00110001000111110110110110010001010", "00110011010011101000100000110001000", "00110101100101100111110111110011100", 
"00110111111110000110101001111110110", "00111010011101010111010100111111010", "00111101000011101101001001101110100", "00111111110001011100010010011011100", 
"01000010100110111001110010101100000", "01000101100100011011100111011011000", "01001000101010011000101111000110100", "01001011111001001001001001101110100", 
"01001111010001000101110110110010000", "01010010110010101001000001100010010", "00000000000000000000000000000000000", "00000000000000000000000000000000000", 
"00000000000000000000000000000000000", "00000000000000000000000000000000000", "00000000000000000000000000000000000", "00000000000000000000000000000000000", 
"00000000000000000000000000000000000", "00000000000000000000000000000000000", "00000000000000000000000000000000000", "00000000000000000000000000000000000", 
"00000000000000000000000000000000000", "00000000000000000000000000000000000", "00000000000000000000000000000000000", "00000000000000000000000000000000000", 
"00000000000000000000000000000000000", "00000000000000000000000000000000000", "00000000000000000000000000000000000", "00000000000000000000000000000000000", 
"00000000000000000000000000000000000", "00000000000000000000000000000000000", "00000000000000000000000000000000000", "00000000000000000000000000000000000", 
"00000000000000000000000000000000000", "00000000000000000000000000000000000", "00000000000000000000000000000000000", "00000000000000000000000000000000000"
);
type calo_calo_cos_dphi_lut_sfixed_array is array (0 to 2**MAX_CALO_PHI_BITS-1) of sfixed(1 downto -20);
constant CALO_CALO_COS_DPHI_LUT_SFIXED : calo_calo_cos_dphi_lut_sfixed_array := (
"0100000000000000000000", "0011111111101111100110", "0011111110111110011100", "0011111101101100100010", 
"0011111100001010001110", "0011111001110110110010", "0011110111010010111100", "0011110100001110010100", 
"0011110000101000111100", "0011101100100010110100", "0011100111111011111000", "0011100011000100100110", 
"0011011101101100100010", "0011010111110011101100", "0011010001101010011110", "0011001011000000100000", 
"0011000100000110001000", "0010111100101011000000", "0010110100111111011110", "0010101101000011100100", 
"0010100100100110111010", "0010011011111001110110", "0010010010111100011010", "0010001001011110001100", 
"0001111111111111111110", "0001110110010001011010", "0001101100010010011010", "0001100010000011000100", 
"0001010111100011010100", "0001001101000011100100", "0001000010010011011100", "0000110111010010111100", 
"0000101100100010110100", "0000100001100010010010", "0000010110010001011010", "0000001011010000111000", 
"0000000000000000000000", "1000001011010000111000", "1000010110010001011010", "1000100001100010010010", 
"1000101100100010110100", "1000110111010010111100", "1001000010010011011100", "1001001101000011100100", 
"1001010111100011010100", "1001100010000011000100", "1001101100010010011010", "1001110110010001011010", 
"1001111111111111111110", "1010001001011110001100", "1010010010111100011010", "1010011011111001110110", 
"1010100100100110111010", "1010101101000011100100", "1010110100111111011110", "1010111100101011000000", 
"1011000100000110001000", "1011001011000000100000", "1011010001101010011110", "1011010111110011101100", 
"1011011101101100100010", "1011100011000100100110", "1011100111111011111000", "1011101100100010110100", 
"1011110000101000111100", "1011110100001110010100", "1011110111010010111100", "1011111001110110110010", 
"1011111100001010001110", "1011111101101100100010", "1011111110111110011100", "1011111111101111100110", 
"1100000000000000000000", "1011111111101111100110", "1011111110111110011100", "1011111101101100100010", 
"1011111100001010001110", "1011111001110110110010", "1011110111010010111100", "1011110100001110010100", 
"1011110000101000111100", "1011101100100010110100", "1011100111111011111000", "1011100011000100100110", 
"1011011101101100100010", "1011010111110011101100", "1011010001101010011110", "1011001011000000100000", 
"1011000100000110001000", "1010111100101011000000", "1010110100111111011110", "1010101101000011100100", 
"1010100100100110111010", "1010011011111001110110", "1010010010111100011010", "1010001001011110001100", 
"1001111111111111111110", "1001110110010001011010", "1001101100010010011010", "1001100010000011000100", 
"1001010111100011010100", "1001001101000011100100", "1001000010010011011100", "1000110111010010111100", 
"1000101100100010110100", "1000100001100010010010", "1000010110010001011010", "1000001011010000111000", 
"0000000000000000000000", "0000001011010000111000", "0000010110010001011010", "0000100001100010010010", 
"0000101100100010110100", "0000110111010010111100", "0001000010010011011100", "0001001101000011100100", 
"0001010111100011010100", "0001100010000011000100", "0001101100010010011010", "0001110110010001011010", 
"0001111111111111111110", "0010001001011110001100", "0010010010111100011010", "0010011011111001110110", 
"0010100100100110111010", "0010101101000011100100", "0010110100111111011110", "0010111100101011000000", 
"0011000100000110001000", "0011001011000000100000", "0011010001101010011110", "0011010111110011101100", 
"0011011101101100100010", "0011100011000100100110", "0011100111111011111000", "0011101100100010110100", 
"0011110000101000111100", "0011110100001110010100", "0011110111010010111100", "0011111001110110110010", 
"0011111100001010001110", "0011111101101100100010", "0011111110111110011100", "0011111111101111100110", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000"
);
type muon_muon_diff_eta_lut_sfixed_array is array (0 to 2**(MUON_ETA_HIGH-MUON_ETA_LOW+1)-1) of sfixed(3 downto -20);
constant MU_MU_DIFF_ETA_LUT_SFIXED : muon_muon_diff_eta_lut_sfixed_array := (
"000000000000000000000000", "000000000010110100001110", "000000000101101000011100", "000000001000011100101010", 
"000000001011010000111000", "000000001101110100101110", "000000010000101000111100", "000000010011011101001010", 
"000000010110010001011010", "000000011001000101101000", "000000011011111001110110", "000000011110101110000100", 
"000000100001100010010010", "000000100100000110001000", "000000100110111010010110", "000000101001101110100100", 
"000000101100100010110100", "000000101111010111000010", "000000110010001011010000", "000000110100111111011110", 
"000000110111100011010100", "000000111010010111100010", "000000111101001011110000", "000000111111111111111110", 
"000001000010110100001110", "000001000101101000011100", "000001001000011100101010", "000001001011010000111000", 
"000001001110000101000110", "000001010000101000111100", "000001010011011101001010", "000001010110010001011010", 
"000001011001000101101000", "000001011011111001110110", "000001011110101110000100", "000001100001100010010010", 
"000001100100000110001000", "000001100110111010010110", "000001101001101110100100", "000001101100100010110100", 
"000001101111010111000010", "000001110010001011010000", "000001110100111111011110", "000001110111110011101100", 
"000001111010100111111010", "000001111101001011110000", "000001111111111111111110", "000010000010110100001110", 
"000010000101101000011100", "000010001000011100101010", "000010001011010000111000", "000010001110000101000110", 
"000010010000111001010110", "000010010011011101001010", "000010010110010001011010", "000010011001000101101000", 
"000010011011111001110110", "000010011110101110000100", "000010100001100010010010", "000010100100010110100000", 
"000010100111001010110000", "000010101001101110100100", "000010101100100010110100", "000010101111010111000010", 
"000010110010001011010000", "000010110100111111011110", "000010110111110011101100", "000010111010100111111010", 
"000010111101001011110000", "000010111111111111111110", "000011000010110100001110", "000011000101101000011100", 
"000011001000011100101010", "000011001011010000111000", "000011001110000101000110", "000011010000111001010110", 
"000011010011011101001010", "000011010110010001011010", "000011011001000101101000", "000011011011111001110110", 
"000011011110101110000100", "000011100001100010010010", "000011100100010110100000", "000011100111001010110000", 
"000011101001111110111110", "000011101100100010110100", "000011101111010111000010", "000011110010001011010000", 
"000011110100111111011110", "000011110111110011101100", "000011111010100111111010", "000011111101011100001010", 
"000100000000010000011000", "000100000010110100001110", "000100000101101000011100", "000100001000011100101010", 
"000100001011010000111000", "000100001110000101000110", "000100010000111001010110", "000100010011101101100100", 
"000100010110100001110010", "000100011001000101101000", "000100011011111001110110", "000100011110101110000100", 
"000100100001100010010010", "000100100100010110100000", "000100100111001010110000", "000100101001111110111110", 
"000100101100100010110100", "000100101111010111000010", "000100110010001011010000", "000100110100111111011110", 
"000100110111110011101100", "000100111010100111111010", "000100111101011100001010", "000101000000010000011000", 
"000101000010110100001110", "000101000101101000011100", "000101001000011100101010", "000101001011010000111000", 
"000101001110000101000110", "000101010000111001010110", "000101010011101101100100", "000101010110100001110010", 
"000101011001000101101000", "000101011011111001110110", "000101011110101110000100", "000101100001100010010010", 
"000101100100010110100000", "000101100111001010110000", "000101101001111110111110", "000101101100110011001100", 
"000101101111100111011010", "000101110010001011010000", "000101110100111111011110", "000101110111110011101100", 
"000101111010100111111010", "000101111101011100001010", "000110000000010000011000", "000110000011000100100110", 
"000110000101111000110100", "000110001000011100101010", "000110001011010000111000", "000110001110000101000110", 
"000110010000111001010110", "000110010011101101100100", "000110010110100001110010", "000110011001010110000000", 
"000110011100001010001110", "000110011110101110000100", "000110100001100010010010", "000110100100010110100000", 
"000110100111001010110000", "000110101001111110111110", "000110101100110011001100", "000110101111100111011010", 
"000110110010011011101000", "000110110100111111011110", "000110110111110011101100", "000110111010100111111010", 
"000110111101011100001010", "000111000000010000011000", "000111000011000100100110", "000111000101111000110100", 
"000111001000011100101010", "000111001011010000111000", "000111001110000101000110", "000111010000111001010110", 
"000111010011101101100100", "000111010110100001110010", "000111011001010110000000", "000111011100001010001110", 
"000111011110101110000100", "000111100001100010010010", "000111100100010110100000", "000111100111001010110000", 
"000111101001111110111110", "000111101100110011001100", "000111101111100111011010", "000111110010011011101000", 
"000111110100111111011110", "000111110111110011101100", "000111111010100111111010", "000111111101011100001010", 
"001000000000010000011000", "001000000011000100100110", "001000000101111000110100", "001000001000101101000010", 
"001000001011010000111000", "001000001110000101000110", "001000010000111001010110", "001000010011101101100100", 
"001000010110100001110010", "001000011001010110000000", "001000011100001010001110", "001000011110111110011100", 
"001000100001110010101100", "001000100100010110100000", "001000100111001010110000", "001000101001111110111110", 
"001000101100110011001100", "001000101111100111011010", "001000110010011011101000", "001000110101001111110110", 
"001000110111110011101100", "001000111010100111111010", "001000111101011100001010", "001001000000010000011000", 
"001001000011000100100110", "001001000101111000110100", "001001001000101101000010", "001001001011100001010000", 
"001001001110010101100000", "001001010000111001010110", "001001010011101101100100", "001001010110100001110010", 
"001001011001010110000000", "001001011100001010001110", "001001011110111110011100", "001001100001110010101100", 
"001001100100010110100000", "001001100111001010110000", "001001101001111110111110", "001001101100110011001100", 
"001001101111100111011010", "001001110010011011101000", "001001110101001111110110", "001001111000000100000110", 
"001001111010111000010100", "001001111101011100001010", "001010000000010000011000", "001010000011000100100110", 
"001010000101111000110100", "001010001000101101000010", "001010001011100001010000", "001010001110010101100000", 
"001010010001001001101110", "001010010011101101100100", "001010010110100001110010", "001010011001010110000000", 
"001010011100001010001110", "001010011110111110011100", "001010100001110010101100", "001010100100100110111010", 
"001010100111001010110000", "001010101001111110111110", "001010101100110011001100", "001010101111100111011010", 
"001010110010011011101000", "001010110101001111110110", "001010111000000100000110", "001010111010111000010100", 
"001010111101101100100010", "001011000000010000011000", "001011000011000100100110", "001011000101111000110100", 
"001011001000101101000010", "001011001011100001010000", "001011001110010101100000", "001011010001001001101110", 
"001011010011101101100100", "001011010110100001110010", "001011011001010110000000", "001011011100001010001110", 
"001011011110111110011100", "001011100001110010101100", "001011100100100110111010", "001011100111011011001000", 
"001011101010001111010110", "001011101100110011001100", "001011101111100111011010", "001011110010011011101000", 
"001011110101001111110110", "001011111000000100000110", "001011111010111000010100", "001011111101101100100010", 
"001100000000010000011000", "001100000011000100100110", "001100000101111000110100", "001100001000101101000010", 
"001100001011100001010000", "001100001110010101100000", "001100010001001001101110", "001100010011111101111100", 
"001100010110110010001010", "001100011001010110000000", "001100011100001010001110", "001100011110111110011100", 
"001100100001110010101100", "001100100100100110111010", "001100100111011011001000", "001100101010001111010110", 
"001100101101000011100100", "001100101111100111011010", "001100110010011011101000", "001100110101001111110110", 
"001100111000000100000110", "001100111010111000010100", "001100111101101100100010", "001101000000100000110000", 
"001101000011000100100110", "001101000101111000110100", "001101001000101101000010", "001101001011100001010000", 
"001101001110010101100000", "001101010001001001101110", "001101010011111101111100", "001101010110110010001010", 
"001101011001100110011000", "001101011100001010001110", "001101011110111110011100", "001101100001110010101100", 
"001101100100100110111010", "001101100111011011001000", "001101101010001111010110", "001101101101000011100100", 
"001101101111100111011010", "001101110010011011101000", "001101110101001111110110", "001101111000000100000110", 
"001101111010111000010100", "001101111101101100100010", "001110000000100000110000", "001110000011010100111110", 
"001110000110001001001100", "001110001000101101000010", "001110001011100001010000", "001110001110010101100000", 
"001110010001001001101110", "001110010011111101111100", "001110010110110010001010", "001110011001100110011000", 
"001110011100001010001110", "001110011110111110011100", "001110100001110010101100", "001110100100100110111010", 
"001110100111011011001000", "001110101010001111010110", "001110101101000011100100", "001110101111110111110010", 
"001110110010101100000010", "001110110101001111110110", "001110111000000100000110", "001110111010111000010100", 
"001110111101101100100010", "001111000000100000110000", "001111000011010100111110", "001111000110001001001100", 
"001111001000101101000010", "001111001011100001010000", "001111001110010101100000", "001111010001001001101110", 
"001111010011111101111100", "001111010110110010001010", "001111011001100110011000", "001111011100011010100110", 
"001111011110111110011100", "001111100001110010101100", "001111100100100110111010", "001111100111011011001000", 
"001111101010001111010110", "001111101101000011100100", "001111101111110111110010", "001111110010101100000010", 
"001111110101100000010000", "001111111000000100000110", "001111111010111000010100", "001111111101101100100010", 
"010000000000100000110000", "010000000011010100111110", "010000000110001001001100", "010000001000111101011100", 
"010000001011100001010000", "010000001110010101100000", "010000010001001001101110", "010000010011111101111100", 
"010000010110110010001010", "010000011001100110011000", "010000011100011010100110", "010000011111001110110110", 
"010000100001110010101100", "010000100100100110111010", "010000100111011011001000", "010000101010001111010110", 
"010000101101000011100100", "010000101111110111110010", "010000110010101100000010", "010000110101100000010000", 
"010000111000010100011110", "010000111010111000010100", "010000111101101100100010", "010001000000100000110000", 
"010001000011010100111110", "010001000110001001001100", "010001001000111101011100", "010001001011110001101010", 
"010001001110100101111000", "010001010001001001101110", "010001010011111101111100", "010001010110110010001010", 
"010001011001100110011000", "010001011100011010100110", "010001011111001110110110", "010001100010000011000100", 
"010001100100100110111010", "010001100111011011001000", "010001101010001111010110", "010001101101000011100100", 
"010001101111110111110010", "010001110010101100000010", "010001110101100000010000", "010001111000010100011110", 
"010001111010111000010100", "010001111101101100100010", "010010000000100000110000", "010010000011010100111110", 
"010010000110001001001100", "010010001000111101011100", "010010001011110001101010", "010010001110100101111000", 
"010010010001011010000110", "010010010011111101111100", "010010010110110010001010", "010010011001100110011000", 
"010010011100011010100110", "010010011111001110110110", "010010100010000011000100", "010010100100110111010010", 
"010010100111101011100000", "010010101010001111010110", "010010101101000011100100", "010010101111110111110010", 
"010010110010101100000010", "010010110101100000010000", "010010111000010100011110", "010010111011001000101100", 
"010010111101101100100010", "010011000000100000110000", "010011000011010100111110", "010011000110001001001100", 
"010011001000111101011100", "010011001011110001101010", "010011001110100101111000", "010011010001011010000110", 
"010011010100001110010100", "010011010110110010001010", "010011011001100110011000", "010011011100011010100110", 
"010011011111001110110110", "010011100010000011000100", "010011100100110111010010", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000"
);
type muon_muon_diff_phi_lut_sfixed_array is array (0 to 2**(MUON_PHI_HIGH-MUON_PHI_LOW+1)-1) of sfixed(3 downto -20);
constant MU_MU_DIFF_PHI_LUT_SFIXED : muon_muon_diff_phi_lut_sfixed_array := (
"000000000000000000000000", "000000000010110100001110", "000000000101101000011100", "000000001000011100101010", 
"000000001011010000111000", "000000001110000101000110", "000000010000101000111100", "000000010011011101001010", 
"000000010110010001011010", "000000011001000101101000", "000000011011111001110110", "000000011110101110000100", 
"000000100001100010010010", "000000100100010110100000", "000000100111001010110000", "000000101001111110111110", 
"000000101100110011001100", "000000101111010111000010", "000000110010001011010000", "000000110100111111011110", 
"000000110111110011101100", "000000111010100111111010", "000000111101011100001010", "000001000000010000011000", 
"000001000011000100100110", "000001000101111000110100", "000001001000101101000010", "000001001011100001010000", 
"000001001110000101000110", "000001010000111001010110", "000001010011101101100100", "000001010110100001110010", 
"000001011001010110000000", "000001011100001010001110", "000001011110111110011100", "000001100001110010101100", 
"000001100100100110111010", "000001100111011011001000", "000001101010001111010110", "000001101100110011001100", 
"000001101111100111011010", "000001110010011011101000", "000001110101001111110110", "000001111000000100000110", 
"000001111010111000010100", "000001111101101100100010", "000010000000100000110000", "000010000011010100111110", 
"000010000110001001001100", "000010001000111101011100", "000010001011100001010000", "000010001110010101100000", 
"000010010001001001101110", "000010010011111101111100", "000010010110110010001010", "000010011001100110011000", 
"000010011100011010100110", "000010011111001110110110", "000010100010000011000100", "000010100100110111010010", 
"000010100111011011001000", "000010101010001111010110", "000010101101000011100100", "000010101111110111110010", 
"000010110010101100000010", "000010110101100000010000", "000010111000010100011110", "000010111011001000101100", 
"000010111101111100111010", "000011000000110001001000", "000011000011100101011000", "000011000110001001001100", 
"000011001000111101011100", "000011001011110001101010", "000011001110100101111000", "000011010001011010000110", 
"000011010100001110010100", "000011010111000010100010", "000011011001110110110010", "000011011100101011000000", 
"000011011111011111001110", "000011100010010011011100", "000011100100110111010010", "000011100111101011100000", 
"000011101010011111101110", "000011101101010011111100", "000011110000001000001100", "000011110010111100011010", 
"000011110101110000101000", "000011111000100100110110", "000011111011011001000100", "000011111110001101010010", 
"000100000001000001100010", "000100000011100101011000", "000100000110011001100110", "000100001001001101110100", 
"000100001100000010000010", "000100001110110110010000", "000100010001101010011110", "000100010100011110101110", 
"000100010111010010111100", "000100011010000111001010", "000100011100111011011000", "000100011111101111100110", 
"000100100010010011011100", "000100100101000111101010", "000100100111111011111000", "000100101010110000001000", 
"000100101101100100010110", "000100110000011000100100", "000100110011001100110010", "000100110110000001000000", 
"000100111000110101001110", "000100111011101001011110", "000100111110011101101100", "000101000001000001100010", 
"000101000011110101110000", "000101000110101001111110", "000101001001011110001100", "000101001100010010011010", 
"000101001111000110101000", "000101010001111010111000", "000101010100101111000110", "000101010111100011010100", 
"000101011010010111100010", "000101011101001011110000", "000101011111101111100110", "000101100010100011110100", 
"000101100101011000000100", "000101101000001100010010", "000101101011000000100000", "000101101101110100101110", 
"000101110000101000111100", "000101110011011101001010", "000101110110010001011010", "000101111001000101101000", 
"000101111011111001110110", "000101111110011101101100", "000110000001010001111010", "000110000100000110001000", 
"000110000110111010010110", "000110001001101110100100", "000110001100100010110100", "000110001111010111000010", 
"000110010010001011010000", "000110010100111111011110", "000110010111110011101100", "000110011010100111111010", 
"000110011101001011110000", "000110011111111111111110", "000110100010110100001110", "000110100101101000011100", 
"000110101000011100101010", "000110101011010000111000", "000110101110000101000110", "000110110000111001010110", 
"000110110011101101100100", "000110110110100001110010", "000110111001010110000000", "000110111011111001110110", 
"000110111110101110000100", "000111000001100010010010", "000111000100010110100000", "000111000111001010110000", 
"000111001001111110111110", "000111001100110011001100", "000111001111100111011010", "000111010010011011101000", 
"000111010101001111110110", "000111011000000100000110", "000111011010100111111010", "000111011101011100001010", 
"000111100000010000011000", "000111100011000100100110", "000111100101111000110100", "000111101000101101000010", 
"000111101011100001010000", "000111101110010101100000", "000111110001001001101110", "000111110011111101111100", 
"000111110110100001110010", "000111111001010110000000", "000111111100001010001110", "000111111110111110011100", 
"001000000001110010101100", "001000000100100110111010", "001000000111011011001000", "001000001010001111010110", 
"001000001101000011100100", "001000001111110111110010", "001000010010101100000010", "001000010101001111110110", 
"001000011000000100000110", "001000011010111000010100", "001000011101101100100010", "001000100000100000110000", 
"001000100011010100111110", "001000100110001001001100", "001000101000111101011100", "001000101011110001101010", 
"001000101110100101111000", "001000110001011010000110", "001000110011111101111100", "001000110110110010001010", 
"001000111001100110011000", "001000111100011010100110", "001000111111001110110110", "001001000010000011000100", 
"001001000100110111010010", "001001000111101011100000", "001001001010011111101110", "001001001101010011111100", 
"001001010000001000001100", "001001010010101100000010", "001001010101100000010000", "001001011000010100011110", 
"001001011011001000101100", "001001011101111100111010", "001001100000110001001000", "001001100011100101011000", 
"001001100110011001100110", "001001101001001101110100", "001001101100000010000010", "001001101110110110010000", 
"001001110001011010000110", "001001110100001110010100", "001001110111000010100010", "001001111001110110110010", 
"001001111100101011000000", "001001111111011111001110", "001010000010010011011100", "001010000101000111101010", 
"001010000111111011111000", "001010001010110000001000", "001010001101100100010110", "001010010000001000001100", 
"001010010010111100011010", "001010010101110000101000", "001010011000100100110110", "001010011011011001000100", 
"001010011110001101010010", "001010100001000001100010", "001010100011110101110000", "001010100110101001111110", 
"001010101001011110001100", "001010101100010010011010", "001010101110110110010000", "001010110001101010011110", 
"001010110100011110101110", "001010110111010010111100", "001010111010000111001010", "001010111100111011011000", 
"001010111111101111100110", "001011000010100011110100", "001011000101011000000100", "001011001000001100010010", 
"001011001011000000100000", "001011001101100100010110", "001011010000011000100100", "001011010011001100110010", 
"001011010110000001000000", "001011011000110101001110", "001011011011101001011110", "001011011110011101101100", 
"001011100001010001111010", "001011100100000110001000", "001011100110111010010110", "001011101001101110100100", 
"001011101100010010011010", "001011101111000110101000", "001011110001111010111000", "001011110100101111000110", 
"001011110111100011010100", "001011111010010111100010", "001011111101001011110000", "001100000000000000000000", 
"001100000010110100001110", "001100000101101000011100", "001100001000011100101010", "001100001011000000100000", 
"001100001101110100101110", "001100010000101000111100", "001100010011011101001010", "001100010110010001011010", 
"001100011001000101101000", "001100011011111001110110", "001100011110101110000100", "001100100001100010010010", 
"001100100100010110100000", "001100100111001010110000", "001100101001101110100100", "001100101100100010110100", 
"001100101111010111000010", "001100110010001011010000", "001100110100111111011110", "001100110111110011101100", 
"001100111010100111111010", "001100111101011100001010", "001101000000010000011000", "001101000011000100100110", 
"001101000101101000011100", "001101001000011100101010", "001101001011010000111000", "001101001110000101000110", 
"001101010000111001010110", "001101010011101101100100", "001101010110100001110010", "001101011001010110000000", 
"001101011100001010001110", "001101011110111110011100", "001101100001110010101100", "001101100100010110100000", 
"001101100111001010110000", "001101101001111110111110", "001101101100110011001100", "001101101111100111011010", 
"001101110010011011101000", "001101110101001111110110", "001101111000000100000110", "001101111010111000010100", 
"001101111101101100100010", "001110000000100000110000", "001110000011000100100110", "001110000101111000110100", 
"001110001000101101000010", "001110001011100001010000", "001110001110010101100000", "001110010001001001101110", 
"001110010011111101111100", "001110010110110010001010", "001110011001100110011000", "001110011100011010100110", 
"001110011111001110110110", "001110100001110010101100", "001110100100100110111010", "001110100111011011001000", 
"001110101010001111010110", "001110101101000011100100", "001110101111110111110010", "001110110010101100000010", 
"001110110101100000010000", "001110111000010100011110", "001110111011001000101100", "001110111101111100111010", 
"001111000000100000110000", "001111000011010100111110", "001111000110001001001100", "001111001000111101011100", 
"001111001011110001101010", "001111001110100101111000", "001111010001011010000110", "001111010100001110010100", 
"001111010111000010100010", "001111011001110110110010", "001111011100101011000000", "001111011111001110110110", 
"001111100010000011000100", "001111100100110111010010", "001111100111101011100000", "001111101010011111101110", 
"001111101101010011111100", "001111110000001000001100", "001111110010111100011010", "001111110101110000101000", 
"001111111000100100110110", "001111111011011001000100", "001111111101111100111010", "010000000000110001001000", 
"010000000011100101011000", "010000000110011001100110", "010000001001001101110100", "010000001100000010000010", 
"010000001110110110010000", "010000010001101010011110", "010000010100011110101110", "010000010111010010111100", 
"010000011010000111001010", "010000011100101011000000", "010000011111011111001110", "010000100010010011011100", 
"010000100101000111101010", "010000100111111011111000", "010000101010110000001000", "010000101101100100010110", 
"010000110000011000100100", "010000110011001100110010", "010000110110000001000000", "010000111000110101001110", 
"010000111011011001000100", "010000111110001101010010", "010001000001000001100010", "010001000011110101110000", 
"010001000110101001111110", "010001001001011110001100", "010001001100010010011010", "010001001111000110101000", 
"010001010001111010111000", "010001010100101111000110", "010001010111100011010100", "010001011010000111001010", 
"010001011100111011011000", "010001011111101111100110", "010001100010100011110100", "010001100101011000000100", 
"010001101000001100010010", "010001101011000000100000", "010001101101110100101110", "010001110000101000111100", 
"010001110011011101001010", "010001110110000001000000", "010001111000110101001110", "010001111011101001011110", 
"010001111110011101101100", "010010000001010001111010", "010010000100000110001000", "010010000110111010010110", 
"010010001001101110100100", "010010001100100010110100", "010010001111010111000010", "010010010010001011010000", 
"010010010100101111000110", "010010010111100011010100", "010010011010010111100010", "010010011101001011110000", 
"010010011111111111111110", "010010100010110100001110", "010010100101101000011100", "010010101000011100101010", 
"010010101011010000111000", "010010101110000101000110", "010010110000111001010110", "010010110011011101001010", 
"010010110110010001011010", "010010111001000101101000", "010010111011111001110110", "010010111110101110000100", 
"010011000001100010010010", "010011000100010110100000", "010011000111001010110000", "010011001001111110111110", 
"010011001100110011001100", "010011001111100111011010", "010011010010001011010000", "010011010100111111011110", 
"010011010111110011101100", "010011011010100111111010", "010011011101011100001010", "010011100000010000011000", 
"010011100011000100100110", "010011100101111000110100", "010011101000101101000010", "010011101011100001010000", 
"010011101110010101100000", "010011110000111001010110", "010011110011101101100100", "010011110110100001110010", 
"010011111001010110000000", "010011111100001010001110", "010011111110111110011100", "010100000001110010101100", 
"010100000100100110111010", "010100000111011011001000", "010100001010001111010110", "010100001101000011100100", 
"010100001111100111011010", "010100010010011011101000", "010100010101001111110110", "010100011000000100000110", 
"010100011010111000010100", "010100011101101100100010", "010100100000100000110000", "010100100011010100111110", 
"010100100110001001001100", "010100101000111101011100", "010100101011110001101010", "010100101110010101100000", 
"010100110001001001101110", "010100110011111101111100", "010100110110110010001010", "010100111001100110011000", 
"010100111100011010100110", "010100111111001110110110", "010101000010000011000100", "010101000100110111010010", 
"010101000111101011100000", "010101001010011111101110", "010101001101000011100100", "010101001111110111110010", 
"010101010010101100000010", "010101010101100000010000", "010101011000010100011110", "010101011011001000101100", 
"010101011101111100111010", "010101100000110001001000", "010101100011100101011000", "010101100110011001100110", 
"010101101001001101110100", "010101101011110001101010", "010101101110100101111000", "010101110001011010000110", 
"010101110100001110010100", "010101110111000010100010", "010101111001110110110010", "010101111100101011000000", 
"010101111111011111001110", "010110000010010011011100", "010110000101000111101010", "010110000111111011111000", 
"010110001010011111101110", "010110001101010011111100", "010110010000001000001100", "010110010010111100011010", 
"010110010101110000101000", "010110011000100100110110", "010110011011011001000100", "010110011110001101010010", 
"010110100001000001100010", "010110100011110101110000", "010110100110101001111110", "010110101001001101110100", 
"010110101100000010000010", "010110101110110110010000", "010110110001101010011110", "010110110100011110101110", 
"010110110111010010111100", "010110111010000111001010", "010110111100111011011000", "010110111111101111100110", 
"010111000010100011110100", "010111000101000111101010", "010111000111111011111000", "010111001010110000001000", 
"010111001101100100010110", "010111010000011000100100", "010111010011001100110010", "010111010110000001000000", 
"010111011000110101001110", "010111011011101001011110", "010111011110011101101100", "010111100001010001111010", 
"010111100011110101110000", "010111100110101001111110", "010111101001011110001100", "010111101100010010011010", 
"010111101111000110101000", "010111110001111010111000", "010111110100101111000110", "010111110111100011010100", 
"010111111010010111100010", "010111111101001011110000", "011000000000000000000000", "011000000010100011110100", 
"011000000101011000000100", "011000001000001100010010", "011000001011000000100000", "011000001101110100101110", 
"011000010000101000111100", "011000010011011101001010", "011000010110010001011010", "011000011001000101101000", 
"011000011011111001110110", "011000011110101110000100", "011000100001010001111010", "011000100100000110001000", 
"011000100110111010010110", "011000101001101110100100", "011000101100100010110100", "011000101111010111000010", 
"011000110010001011010000", "011000110100111111011110", "011000110111110011101100", "011000111010100111111010", 
"011000111101011100001010", "011000111111111111111110", "011001000010110100001110", "011001000101101000011100", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000", 
"000000000000000000000000", "000000000000000000000000", "000000000000000000000000", "000000000000000000000000"
);
type muon_muon_cosh_deta_lut_sfixed_array is array (0 to 2**(MUON_ETA_HIGH-MUON_ETA_LOW+1)-1) of sfixed(7 downto -20);
constant MU_MU_COSH_DETA_LUT_SFIXED : muon_muon_cosh_deta_lut_sfixed_array := (
"0000000100000000000000000000", "0000000100000000000001101000", "0000000100000000000011010000", "0000000100000000001000001100", 
"0000000100000000001110101110", "0000000100000000011000100100", "0000000100000000100010011010", "0000000100000000101111100000", 
"0000000100000000111110010000", "0000000100000001001110101000", "0000000100000001100000101010", "0000000100000001110101111100", 
"0000000100000010001011010000", "0000000100000010100011110100", "0000000100000010111110000010", "0000000100000011011001111010", 
"0000000100000011111001000010", "0000000100000100011000001010", "0000000100000100111010100100", "0000000100000101011110100110", 
"0000000100000110000100010010", "0000000100000110101101010000", "0000000100000111010111110110", "0000000100001000000010011100", 
"0000000100001000110001111110", "0000000100001001100001011110", "0000000100001010010010101000", "0000000100001011000111000100", 
"0000000100001011111101001000", "0000000100001100110100110100", "0000000100001101101111110100", "0000000100001110101100011100", 
"0000000100001111101010101100", "0000000100010000101010100110", "0000000100010001101100001000", "0000000100010010110000111100", 
"0000000100010011110111011000", "0000000100010101000001001000", "0000000100010110001010110110", "0000000100010111010111110110", 
"0000000100011000100110100000", "0000000100011001111000011010", "0000000100011011001010010100", "0000000100011100011111100010", 
"0000000100011101111000000000", "0000000100011111010010000110", "0000000100100000101101111000", "0000000100100010001011010000", 
"0000000100100011101011111010", "0000000100100101001110001110", "0000000100100110110010001010", "0000000100101000011001011000", 
"0000000100101010000010010000", "0000000100101011101110011000", "0000000100101101011010100000", "0000000100101111001011100100", 
"0000000100110000111100100110", "0000000100110010110010100100", "0000000100110100101000100010", "0000000100110110100001110010", 
"0000000100111000011100101010", "0000000100111010011010110100", "0000000100111100011010100110", "0000000100111110011101101100", 
"0000000101000000100010011010", "0000000101000010101010011000", "0000000101000100110100000000", "0000000101000111000000111010", 
"0000000101001001001111011100", "0000000101001011100001010000", "0000000101001101110100101110", "0000000101010000001011011110", 
"0000000101010010100011110100", "0000000101010100111111011110", "0000000101010111011110011010", "0000000101011001111110111110", 
"0000000101011100100001001010", "0000000101011111001000010010", "0000000101100001110001000010", "0000000101100100011011011100", 
"0000000101100111001001000110", "0000000101101001111010000010", "0000000101101100101110010010", "0000000101101111100100001000", 
"0000000101110010011101010010", "0000000101110101011000000100", "0000000101111000010111110000", "0000000101111011011001000100", 
"0000000101111110011101101100", "0000000110000001100011111100", "0000000110000100101111000110", "0000000110000111111011111000", 
"0000000110001011001011111110", "0000000110001110011101101100", "0000000110010001110100010100", "0000000110010101001110001110", 
"0000000110011000101001110000", "0000000110011100001000100110", "0000000110011111101010101100", "0000000110100011010001101100", 
"0000000110100110111010010110", "0000000110101010100110010010", "0000000110101110010011110110", "0000000110110010000110010110", 
"0000000110110101111100000110", "0000000110111001110101001000", "0000000110111101110001011100", "0000000111000001110001000010", 
"0000000111000101110011111010", "0000000111001001111011101100", "0000000111001110000101000110", "0000000111010010010011011100", 
"0000000111010110100011011010", "0000000111011010111000010100", "0000000111011111010000011110", "0000000111100011101011111010", 
"0000000111101000001100010010", "0000000111101100101110010010", "0000000111110001010101001100", "0000000111110110000001000000", 
"0000000111111010101110011110", "0000000111111111100000110110", "0000001000000100011000001010", "0000001000001001010001000110", 
"0000001000001110001110111100", "0000001000010011010001101100", "0000001000011000010111110000", "0000001000011101100001000100", 
"0000001000100010101111010010", "0000001000101000000010011100", "0000001000101101011000111000", "0000001000110010110010100100", 
"0000001000111000010010110100", "0000001000111101110110010110", "0000001001000011011101001010", "0000001001001001001000111010", 
"0000001001001110111001100010", "0000001001010100101111000110", "0000001001011010100111111010", "0000001001100000100101101010", 
"0000001001100110101000010110", "0000001001101100101111111010", "0000001001110010111100011010", "0000001001111001001100001010", 
"0000001001111111100010100000", "0000001010000101111100000110", "0000001010001100011100010000", "0000001010010010111111101100", 
"0000001010011001101000000010", "0000001010100000010110111100", "0000001010100111001010110000", "0000001010101110000011011110", 
"0000001010110100111111011110", "0000001010111100000011101010", "0000001011000011001011001010", "0000001011001010011001001100", 
"0000001011010001101100001000", "0000001011011001000011111110", "0000001011100000100010011010", "0000001011101000000101101110", 
"0000001011101111101101111110", "0000001011110111011100110000", "0000001011111111010010000110", "0000001100000111001100011000", 
"0000001100001111001011100100", "0000001100010111010010111100", "0000001100011111011111001110", "0000001100100111110000011010", 
"0000001100110000001001110100", "0000001100111000101000001000", "0000001101000001001101000000", "0000001101001001110110110010", 
"0000001101010010101000110000", "0000001101011011100001010000", "0000001101100100011110101110", "0000001101101101100100010110", 
"0000001101110110101110111000", "0000001110000000000001101000", "0000001110001001011010111010", "0000001110010010111010110000", 
"0000001110011100100001001010", "0000001110100110001111110000", "0000001110110000000011010000", "0000001110111010000000100110", 
"0000001111000100000010110110", "0000001111001110001101010010", "0000001111011000011111111100", "0000001111100010111001001000", 
"0000001111101101011010100000", "0000001111111000000010011100", "0000010000000010110010100100", "0000010000001101101010111000", 
"0000010000011000101001110000", "0000010000100011110010011110", "0000010000101111000001101110", "0000010000111010011010110100", 
"0000010001000101111010011110", "0000010001010001100010010010", "0000010001011101010011111100", "0000010001101001001100001010", 
"0000010001110101001110001110", "0000010010000001011000011110", "0000010010001101101010111000", "0000010010011010000111001010", 
"0000010010100110101101010000", "0000010010110011011001111010", "0000010011000000010010000000", "0000010011001101010000101100", 
"0000010011011010011010110100", "0000010011100111101101001010", "0000010011110101001010111100", "0000010100000010110000111100", 
"0000010100010000100000110000", "0000010100011110011000110000", "0000010100101100011100010000", "0000010100111010101001100100", 
"0000010101001001000010010110", "0000010101010111100011010100", "0000010101100110001111110000", "0000010101110101000110000010", 
"0000010110000100000111110010", "0000010110010011010011010110", "0000010110100010101010011000", "0000010110110010001100111000", 
"0000010111000001111001001110", "0000010111010001110001000010", "0000010111100001110100010100", "0000010111110010000011000100", 
"0000011000000010011011101000", "0000011000010011000001010100", "0000011000100011110100000110", "0000011000110100110000101110", 
"0000011001000101111010011110", "0000011001010111001111101010", "0000011001101000110001111110", "0000011001111010011111101110", 
"0000011010001100011010100110", "0000011010011110100010100110", "0000011010110000110110000100", "0000011011000011011000010000", 
"0000011011010110000101111100", "0000011011101001000000101100", "0000011011111100001010001110", "0000011100001111100000110110", 
"0000011100100011000100100110", "0000011100110110110111000100", "0000011101001010110110101010", "0000011101011111000101000000", 
"0000011101110011100010000110", "0000011110001000001100010010", "0000011110011101000110110110", "0000011110110010001110100010", 
"0000011111000111100100111100", "0000011111011101001011110000", "0000011111110011000001010100", "0000100000001001000101101000", 
"0000100000011111011010010100", "0000100000110101111111011000", "0000100001001100110011001100", "0000100001100011110111011000", 
"0000100001111011001011111110", "0000100010010010101111010010", "0000100010101010100110010010", "0000100011000010101100000010", 
"0000100011011011000011110010", "0000100011110011101011111010", "0000100100001100100100011100", "0000100100100101110000101000", 
"0000100100111111001101001100", "0000100101011000111011110010", "0000100101110010111110000010", "0000100110001101010000101100", 
"0000100110100111110110111110", "0000100111000010101111010010", "0000100111011101111011010010", "0000100111111001011001010010", 
"0000101000010101001010111100", "0000101000110001010000010010", "0000101001001101101001010000", "0000101001101010010111100010", 
"0000101010000111010111110110", "0000101010100100101101011100", "0000101011000010011000010110", "0000101011100000010110111100", 
"0000101011111110101100011100", "0000101100011101010101100110", "0000101100111100010100000100", "0000101101011011101001011110", 
"0000101101111011010100001010", "0000101110011011010101110010", "0000101110111011101100101110", "0000101111011100011010100110", 
"0000101111111101100001000100", "0000110000011110111100110100", "0000110001000000110001001000", "0000110001100010111110000010", 
"0000110010000101100000010000", "0000110010101000011100101010", "0000110011001011110001101010", "0000110011101111011111001110", 
"0000110100010011100101011000", "0000110100111000000101101110", "0000110101011100111110101010", "0000110110000010010001110100", 
"0000110110100111111111001010", "0000110111001110001000011000", "0000110111110100101010001100", "0000111000011011100111110100", 
"0000111001000011000001010100", "0000111001101010110110101010", "0000111010010011000110001110", "0000111010111011110011010010", 
"0000111011100100111100001100", "0000111100001110100010100110", "0000111100111000100110100000", "0000111101100011000111111000", 
"0000111110001110000110110000", "0000111110111001100011000110", "0000111111100101011110100110", "0001000000010001111001001110", 
"0001000000111110110010111110", "0001000001101100001011111000", "0001000010011010000011111000", "0001000011001000011100101010", 
"0001000011110111010110001110", "0001000100100110110000100010", "0001000101010110101011100110", "0001000110000111001001000110", 
"0001000110111000000111010110", "0001000111101001101001101010", "0001001000011011101100101110", "0001001001001110010011110110", 
"0001001010000001011111000000", "0001001010110101001100100110", "0001001011101001011111110110", "0001001100011110010111001000", 
"0001001101010011110100000110", "0001001110001001110101001000", "0001001111000000011101011110", "0001001111110111101011100000", 
"0001010000101111011111001110", "0001010001100111111011111000", "0001010010100000111111111000", "0001010011011010101011001100", 
"0001010100010100111101110110", "0001010101001111111011000100", "0001010110001011100001010000", "0001010111000111110000011010", 
"0001011000000100101010001100", "0001011001000010001110100010", "0001011010000000011101011110", "0001011010111111011000101010", 
"0001011011111111000000000110", "0001011100111111010011110000", "0001011110000000010101010010", "0001011111000010000011000100", 
"0001100000000100100000010110", "0001100001000111101011100000", "0001100010001011100100100010", "0001100011010000001110101110", 
"0001100100010101101000011100", "0001100101011011110011010010", "0001100110100010101101101010", "0001100111101010011010110100", 
"0001101000110010111010110000", "0001101001111100001101100000", "0001101011000110010001011010", "0001101100010001001011010110", 
"0001101101011100111001110000", "0001101110101001011100100100", "0001101111110110110011110100", "0001110001000101000010110000", 
"0001110010010100000111110010", "0001110011100100000100100000", "0001110100110100111000111010", "0001110110000110100110101100", 
"0001110111011001001101110100", "0001111000101100101110010010", "0001111010000001001000000100", "0001111011010110011110100000", 
"0001111100101100101111111010", "0001111110000011111101111100", "0001111111011100001000100110", "0010000000110101010001100000", 
"0010000010001111011000101010", "0010000011101010011111101110", "0010000101000110100101000100", "0010000110100011101011111010", 
"0010001000000001110100010100", "0010001001100000111110010000", "0010001011000001001001101110", "0010001100100010011010000000", 
"0010001110000100101101011100", "0010001111101000000101101110", "0010010001001100100100011100", "0010010010110010000111111110", 
"0010010100011000110011100110", "0010010110000000100111010100", "0010010111101001100011000110", "0010011001010011101000101000", 
"0010011010111110111001100010", "0010011100101011010100001010", "0010011110011000111011110010", "0010100000000111101110110010", 
"0010100001110111110000011010", "0010100011101000111111000100", "0010100101011011011110000000", "0010100111001111001101001100", 
"0010101001000100001100101100", "0010101010111010011110000110", "0010101100110010000011000100", "0010101110101010111011100110", 
"0010110000100101001001010100", "0010110010100000101010100110", "0010110100011101100100010110", "0010110110011011110100111100", 
"0010111000011011011110000000", "0010111010011100011111100010", "0010111100011110111011001010", "0010111110100010110100001110", 
"0011000000101000000111010110", "0011000010101110111001100010", "0011000100110111001001000110", "0011000111000000110111101100", 
"0011001001001100000110111100", "0011001011011000111000100000", "0011001101100111001010110000", "0011001111110111000010100010", 
"0011010010001000011110010010", "0011010100011011011111101000", "0011010110110000001000001100", "0011011001000110010111111100", 
"0011011011011110010010001110", "0011011101110111110110111110", "0011100000010011000110001110", "0011100010110000000001101000", 
"0011100101001110101100011100", "0011100111101111000101000000", "0011101010010001001110101000", "0011101100110101001001010100", 
"0011101111011010110110101010", "0011110010000010010110101110", "0011110100101011101110011000", "0011110111010110111100000000", 
"0011111010000011111111100100", "0011111100110010111110000010", "0011111111100011110111011000", "0100000010010110101011100110", 
"0100000101001011011100010110", "0100001000000010001100111000", "0100001010111010111101001110", "0000000000000000000000000000", 
"0000000000000000000000000000", "0000000000000000000000000000", "0000000000000000000000000000", "0000000000000000000000000000", 
"0000000000000000000000000000", "0000000000000000000000000000", "0000000000000000000000000000", "0000000000000000000000000000", 
"0000000000000000000000000000", "0000000000000000000000000000", "0000000000000000000000000000", "0000000000000000000000000000", 
"0000000000000000000000000000", "0000000000000000000000000000", "0000000000000000000000000000", "0000000000000000000000000000", 
"0000000000000000000000000000", "0000000000000000000000000000", "0000000000000000000000000000", "0000000000000000000000000000", 
"0000000000000000000000000000", "0000000000000000000000000000", "0000000000000000000000000000", "0000000000000000000000000000", 
"0000000000000000000000000000", "0000000000000000000000000000", "0000000000000000000000000000", "0000000000000000000000000000", 
"0000000000000000000000000000", "0000000000000000000000000000", "0000000000000000000000000000", "0000000000000000000000000000", 
"0000000000000000000000000000", "0000000000000000000000000000", "0000000000000000000000000000", "0000000000000000000000000000", 
"0000000000000000000000000000", "0000000000000000000000000000", "0000000000000000000000000000", "0000000000000000000000000000", 
"0000000000000000000000000000", "0000000000000000000000000000", "0000000000000000000000000000", "0000000000000000000000000000", 
"0000000000000000000000000000", "0000000000000000000000000000", "0000000000000000000000000000", "0000000000000000000000000000", 
"0000000000000000000000000000", "0000000000000000000000000000", "0000000000000000000000000000", "0000000000000000000000000000", 
"0000000000000000000000000000", "0000000000000000000000000000", "0000000000000000000000000000", "0000000000000000000000000000", 
"0000000000000000000000000000", "0000000000000000000000000000", "0000000000000000000000000000", "0000000000000000000000000000"
);
type muon_muon_cos_dphi_lut_sfixed_array is array (0 to 2**(MUON_PHI_HIGH-MUON_PHI_LOW+1)-1) of sfixed(1 downto -20);
constant MU_MU_COS_DPHI_LUT_SFIXED : muon_muon_cos_dphi_lut_sfixed_array := (
"0100000000000000000000", "0011111111111110010110", "0011111111111100101110", "0011111111110111110010", 
"0011111111101111100110", "0011111111100111011010", "0011111111011101100100", "0011111111010000011110", 
"0011111111000001101110", "0011111110110001010110", "0011111110011111010100", "0011111110001010000010", 
"0011111101110011000110", "0011111101011100001010", "0011111101000001111100", "0011111100100100011100", 
"0011111100000110111100", "0011111011100111110100", "0011111011000101011010", "0011111010100001011000", 
"0011111001111011101100", "0011111001010100011000", "0011111000101001110000", "0011110111111111001010", 
"0011110111010001010010", "0011110110100001110010", "0011110101110000101000", "0011110100111101110110", 
"0011110100001001011010", "0011110011010011010110", "0011110010011010000000", "0011110001100000101010", 
"0011110000100100000010", "0011101111100101110010", "0011101110100101111000", "0011101101100100010110", 
"0011101100100001001010", "0011101011011100010110", "0011101010010100010000", "0011101001001100001010", 
"0011101000000000110100", "0011100110110011110100", "0011100101100110110010", "0011100100010110100000", 
"0011100011000100100110", "0011100001110001000010", "0011100000011011110110", "0011011111000101000000", 
"0011011101101100100010", "0011011100010010011010", "0011011010110110101010", "0011011001011001010010", 
"0011010111111010010000", "0011010110011001100110", "0011010100110111010010", "0011010011010011010110", 
"0011010001101101110000", "0011010000000100111010", "0011001110011100000010", "0011001100110001100010", 
"0011001011000111000100", "0011001001011001010010", "0011000111101001111000", "0011000101111000110100", 
"0011000100000110001000", "0011000010010011011100", "0011000000011101011110", "0010111110100111100000", 
"0010111100101111111010", "0010111010110110101010", "0010111000111011110010", "0010110110111111010010", 
"0010110101000001001000", "0010110011000010111110", "0010110001000001100010", "0010101111000000000110", 
"0010101100111101000000", "0010101010111000010100", "0010101000110001111110", "0010100110101011100110", 
"0010100100100011101000", "0010100010011010000000", "0010100000001110101110", "0010011110000011011110", 
"0010011011110110100100", "0010011001101000000010", "0010010111010111110110", "0010010101000111101010", 
"0010010010110101110110", "0010010000100010011010", "0010001110001110111100", "0010001011111001110110", 
"0010001001100011000110", "0010000111001100011000", "0010000100110100000000", "0010000010011010000000", 
"0001111111111111111110", "0001111101100100010110", "0001111011001000101100", "0001111000101011011010", 
"0001110110001100011110", "0001110011101101100100", "0001110001001110101000", "0001101110101110000100", 
"0001101100001011111000", "0001101001101001101010", "0001100111000101110100", "0001100100100001111110", 
"0001100001111110001010", "0001011111011000101010", "0001011100110001100010", "0001011010001100000100", 
"0001010111100011010100", "0001010100111010100100", "0001010010010001110100", "0001001111101001000010", 
"0001001100111110101010", "0001001010010100010000", "0001000111101000001110", "0001000100111100001100", 
"0001000010010000001010", "0000111111100100001000", "0000111100110110011110", "0000111010001000110010", 
"0000110111011001011110", "0000110100101011110100", "0000110001111100100000", "0000101111001101001100", 
"0000101100011100010000", "0000101001101100111100", "0000100110111100000000", "0000100100001011000010", 
"0000100001011010000110", "0000011110101001001010", "0000011011111000001100", "0000011001000101101000", 
"0000010110010100101010", "0000010011100010000110", "0000010000101111100000", "0000001101111100111010", 
"0000001011001010010100", "0000001000010111110000", "0000000101100101001010", "0000000010110010100100", 
"0000000000000000000000", "1000000010110010100100", "1000000101100101001010", "1000001000010111110000", 
"1000001011001010010100", "1000001101111100111010", "1000010000101111100000", "1000010011100010000110", 
"1000010110010100101010", "1000011001000101101000", "1000011011111000001100", "1000011110101001001010", 
"1000100001011010000110", "1000100100001011000010", "1000100110111100000000", "1000101001101100111100", 
"1000101100011100010000", "1000101111001101001100", "1000110001111100100000", "1000110100101011110100", 
"1000110111011001011110", "1000111010001000110010", "1000111100110110011110", "1000111111100100001000", 
"1001000010010000001010", "1001000100111100001100", "1001000111101000001110", "1001001010010100010000", 
"1001001100111110101010", "1001001111101001000010", "1001010010010001110100", "1001010100111010100100", 
"1001010111100011010100", "1001011010001100000100", "1001011100110001100010", "1001011111011000101010", 
"1001100001111110001010", "1001100100100001111110", "1001100111000101110100", "1001101001101001101010", 
"1001101100001011111000", "1001101110101110000100", "1001110001001110101000", "1001110011101101100100", 
"1001110110001100011110", "1001111000101011011010", "1001111011001000101100", "1001111101100100010110", 
"1001111111111111111110", "1010000010011010000000", "1010000100110100000000", "1010000111001100011000", 
"1010001001100011000110", "1010001011111001110110", "1010001110001110111100", "1010010000100010011010", 
"1010010010110101110110", "1010010101000111101010", "1010010111010111110110", "1010011001101000000010", 
"1010011011110110100100", "1010011110000011011110", "1010100000001110101110", "1010100010011010000000", 
"1010100100100011101000", "1010100110101011100110", "1010101000110001111110", "1010101010111000010100", 
"1010101100111101000000", "1010101111000000000110", "1010110001000001100010", "1010110011000010111110", 
"1010110101000001001000", "1010110110111111010010", "1010111000111011110010", "1010111010110110101010", 
"1010111100101111111010", "1010111110100111100000", "1011000000011101011110", "1011000010010011011100", 
"1011000100000110001000", "1011000101111000110100", "1011000111101001111000", "1011001001011001010010", 
"1011001011000111000100", "1011001100110001100010", "1011001110011100000010", "1011010000000100111010", 
"1011010001101101110000", "1011010011010011010110", "1011010100110111010010", "1011010110011001100110", 
"1011010111111010010000", "1011011001011001010010", "1011011010110110101010", "1011011100010010011010", 
"1011011101101100100010", "1011011111000101000000", "1011100000011011110110", "1011100001110001000010", 
"1011100011000100100110", "1011100100010110100000", "1011100101100110110010", "1011100110110011110100", 
"1011101000000000110100", "1011101001001100001010", "1011101010010100010000", "1011101011011100010110", 
"1011101100100001001010", "1011101101100100010110", "1011101110100101111000", "1011101111100101110010", 
"1011110000100100000010", "1011110001100000101010", "1011110010011010000000", "1011110011010011010110", 
"1011110100001001011010", "1011110100111101110110", "1011110101110000101000", "1011110110100001110010", 
"1011110111010001010010", "1011110111111111001010", "1011111000101001110000", "1011111001010100011000", 
"1011111001111011101100", "1011111010100001011000", "1011111011000101011010", "1011111011100111110100", 
"1011111100000110111100", "1011111100100100011100", "1011111101000001111100", "1011111101011100001010", 
"1011111101110011000110", "1011111110001010000010", "1011111110011111010100", "1011111110110001010110", 
"1011111111000001101110", "1011111111010000011110", "1011111111011101100100", "1011111111100111011010", 
"1011111111101111100110", "1011111111110111110010", "1011111111111100101110", "1011111111111110010110", 
"1100000000000000000000", "1011111111111110010110", "1011111111111100101110", "1011111111110111110010", 
"1011111111101111100110", "1011111111100111011010", "1011111111011101100100", "1011111111010000011110", 
"1011111111000001101110", "1011111110110001010110", "1011111110011111010100", "1011111110001010000010", 
"1011111101110011000110", "1011111101011100001010", "1011111101000001111100", "1011111100100100011100", 
"1011111100000110111100", "1011111011100111110100", "1011111011000101011010", "1011111010100001011000", 
"1011111001111011101100", "1011111001010100011000", "1011111000101001110000", "1011110111111111001010", 
"1011110111010001010010", "1011110110100001110010", "1011110101110000101000", "1011110100111101110110", 
"1011110100001001011010", "1011110011010011010110", "1011110010011010000000", "1011110001100000101010", 
"1011110000100100000010", "1011101111100101110010", "1011101110100101111000", "1011101101100100010110", 
"1011101100100001001010", "1011101011011100010110", "1011101010010100010000", "1011101001001100001010", 
"1011101000000000110100", "1011100110110011110100", "1011100101100110110010", "1011100100010110100000", 
"1011100011000100100110", "1011100001110001000010", "1011100000011011110110", "1011011111000101000000", 
"1011011101101100100010", "1011011100010010011010", "1011011010110110101010", "1011011001011001010010", 
"1011010111111010010000", "1011010110011001100110", "1011010100110111010010", "1011010011010011010110", 
"1011010001101101110000", "1011010000000100111010", "1011001110011100000010", "1011001100110001100010", 
"1011001011000111000100", "1011001001011001010010", "1011000111101001111000", "1011000101111000110100", 
"1011000100000110001000", "1011000010010011011100", "1011000000011101011110", "1010111110100111100000", 
"1010111100101111111010", "1010111010110110101010", "1010111000111011110010", "1010110110111111010010", 
"1010110101000001001000", "1010110011000010111110", "1010110001000001100010", "1010101111000000000110", 
"1010101100111101000000", "1010101010111000010100", "1010101000110001111110", "1010100110101011100110", 
"1010100100100011101000", "1010100010011010000000", "1010100000001110101110", "1010011110000011011110", 
"1010011011110110100100", "1010011001101000000010", "1010010111010111110110", "1010010101000111101010", 
"1010010010110101110110", "1010010000100010011010", "1010001110001110111100", "1010001011111001110110", 
"1010001001100011000110", "1010000111001100011000", "1010000100110100000000", "1010000010011010000000", 
"1001111111111111111110", "1001111101100100010110", "1001111011001000101100", "1001111000101011011010", 
"1001110110001100011110", "1001110011101101100100", "1001110001001110101000", "1001101110101110000100", 
"1001101100001011111000", "1001101001101001101010", "1001100111000101110100", "1001100100100001111110", 
"1001100001111110001010", "1001011111011000101010", "1001011100110001100010", "1001011010001100000100", 
"1001010111100011010100", "1001010100111010100100", "1001010010010001110100", "1001001111101001000010", 
"1001001100111110101010", "1001001010010100010000", "1001000111101000001110", "1001000100111100001100", 
"1001000010010000001010", "1000111111100100001000", "1000111100110110011110", "1000111010001000110010", 
"1000110111011001011110", "1000110100101011110100", "1000110001111100100000", "1000101111001101001100", 
"1000101100011100010000", "1000101001101100111100", "1000100110111100000000", "1000100100001011000010", 
"1000100001011010000110", "1000011110101001001010", "1000011011111000001100", "1000011001000101101000", 
"1000010110010100101010", "1000010011100010000110", "1000010000101111100000", "1000001101111100111010", 
"1000001011001010010100", "1000001000010111110000", "1000000101100101001010", "1000000010110010100100", 
"0000000000000000000000", "0000000010110010100100", "0000000101100101001010", "0000001000010111110000", 
"0000001011001010010100", "0000001101111100111010", "0000010000101111100000", "0000010011100010000110", 
"0000010110010100101010", "0000011001000101101000", "0000011011111000001100", "0000011110101001001010", 
"0000100001011010000110", "0000100100001011000010", "0000100110111100000000", "0000101001101100111100", 
"0000101100011100010000", "0000101111001101001100", "0000110001111100100000", "0000110100101011110100", 
"0000110111011001011110", "0000111010001000110010", "0000111100110110011110", "0000111111100100001000", 
"0001000010010000001010", "0001000100111100001100", "0001000111101000001110", "0001001010010100010000", 
"0001001100111110101010", "0001001111101001000010", "0001010010010001110100", "0001010100111010100100", 
"0001010111100011010100", "0001011010001100000100", "0001011100110001100010", "0001011111011000101010", 
"0001100001111110001010", "0001100100100001111110", "0001100111000101110100", "0001101001101001101010", 
"0001101100001011111000", "0001101110101110000100", "0001110001001110101000", "0001110011101101100100", 
"0001110110001100011110", "0001111000101011011010", "0001111011001000101100", "0001111101100100010110", 
"0001111111111111111110", "0010000010011010000000", "0010000100110100000000", "0010000111001100011000", 
"0010001001100011000110", "0010001011111001110110", "0010001110001110111100", "0010010000100010011010", 
"0010010010110101110110", "0010010101000111101010", "0010010111010111110110", "0010011001101000000010", 
"0010011011110110100100", "0010011110000011011110", "0010100000001110101110", "0010100010011010000000", 
"0010100100100011101000", "0010100110101011100110", "0010101000110001111110", "0010101010111000010100", 
"0010101100111101000000", "0010101111000000000110", "0010110001000001100010", "0010110011000010111110", 
"0010110101000001001000", "0010110110111111010010", "0010111000111011110010", "0010111010110110101010", 
"0010111100101111111010", "0010111110100111100000", "0011000000011101011110", "0011000010010011011100", 
"0011000100000110001000", "0011000101111000110100", "0011000111101001111000", "0011001001011001010010", 
"0011001011000111000100", "0011001100110001100010", "0011001110011100000010", "0011010000000100111010", 
"0011010001101101110000", "0011010011010011010110", "0011010100110111010010", "0011010110011001100110", 
"0011010111111010010000", "0011011001011001010010", "0011011010110110101010", "0011011100010010011010", 
"0011011101101100100010", "0011011111000101000000", "0011100000011011110110", "0011100001110001000010", 
"0011100011000100100110", "0011100100010110100000", "0011100101100110110010", "0011100110110011110100", 
"0011101000000000110100", "0011101001001100001010", "0011101010010100010000", "0011101011011100010110", 
"0011101100100001001010", "0011101101100100010110", "0011101110100101111000", "0011101111100101110010", 
"0011110000100100000010", "0011110001100000101010", "0011110010011010000000", "0011110011010011010110", 
"0011110100001001011010", "0011110100111101110110", "0011110101110000101000", "0011110110100001110010", 
"0011110111010001010010", "0011110111111111001010", "0011111000101001110000", "0011111001010100011000", 
"0011111001111011101100", "0011111010100001011000", "0011111011000101011010", "0011111011100111110100", 
"0011111100000110111100", "0011111100100100011100", "0011111101000001111100", "0011111101011100001010", 
"0011111101110011000110", "0011111110001010000010", "0011111110011111010100", "0011111110110001010110", 
"0011111111000001101110", "0011111111010000011110", "0011111111011101100100", "0011111111100111011010", 
"0011111111101111100110", "0011111111110111110010", "0011111111111100101110", "0011111111111110010110", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000", 
"0000000000000000000000", "0000000000000000000000", "0000000000000000000000", "0000000000000000000000"
);
constant EG_EG_DIFF_ETA_LUT_SFIXED : calo_calo_diff_eta_lut_sfixed_array := CALO_CALO_DIFF_ETA_LUT_SFIXED;
constant EG_TAU_DIFF_ETA_LUT_SFIXED : calo_calo_diff_eta_lut_sfixed_array := CALO_CALO_DIFF_ETA_LUT_SFIXED;
constant EG_JET_DIFF_ETA_LUT_SFIXED : calo_calo_diff_eta_lut_sfixed_array := CALO_CALO_DIFF_ETA_LUT_SFIXED;
constant JET_EG_DIFF_ETA_LUT_SFIXED : calo_calo_diff_eta_lut_sfixed_array := CALO_CALO_DIFF_ETA_LUT_SFIXED;
constant JET_JET_DIFF_ETA_LUT_SFIXED : calo_calo_diff_eta_lut_sfixed_array := CALO_CALO_DIFF_ETA_LUT_SFIXED;
constant JET_TAU_DIFF_ETA_LUT_SFIXED : calo_calo_diff_eta_lut_sfixed_array := CALO_CALO_DIFF_ETA_LUT_SFIXED;
constant TAU_EG_DIFF_ETA_LUT_SFIXED : calo_calo_diff_eta_lut_sfixed_array := CALO_CALO_DIFF_ETA_LUT_SFIXED;
constant TAU_JET_DIFF_ETA_LUT_SFIXED : calo_calo_diff_eta_lut_sfixed_array := CALO_CALO_DIFF_ETA_LUT_SFIXED;
constant TAU_TAU_DIFF_ETA_LUT_SFIXED : calo_calo_diff_eta_lut_sfixed_array := CALO_CALO_DIFF_ETA_LUT_SFIXED;
constant EG_EG_DIFF_PHI_LUT_SFIXED : calo_calo_diff_phi_lut_sfixed_array := CALO_CALO_DIFF_PHI_LUT_SFIXED;
constant EG_TAU_DIFF_PHI_LUT_SFIXED : calo_calo_diff_phi_lut_sfixed_array := CALO_CALO_DIFF_PHI_LUT_SFIXED;
constant EG_JET_DIFF_PHI_LUT_SFIXED : calo_calo_diff_phi_lut_sfixed_array := CALO_CALO_DIFF_PHI_LUT_SFIXED;
constant JET_EG_DIFF_PHI_LUT_SFIXED : calo_calo_diff_phi_lut_sfixed_array := CALO_CALO_DIFF_PHI_LUT_SFIXED;
constant JET_JET_DIFF_PHI_LUT_SFIXED : calo_calo_diff_phi_lut_sfixed_array := CALO_CALO_DIFF_PHI_LUT_SFIXED;
constant JET_TAU_DIFF_PHI_LUT_SFIXED : calo_calo_diff_phi_lut_sfixed_array := CALO_CALO_DIFF_PHI_LUT_SFIXED;
constant TAU_EG_DIFF_PHI_LUT_SFIXED : calo_calo_diff_phi_lut_sfixed_array := CALO_CALO_DIFF_PHI_LUT_SFIXED;
constant TAU_JET_DIFF_PHI_LUT_SFIXED : calo_calo_diff_phi_lut_sfixed_array := CALO_CALO_DIFF_PHI_LUT_SFIXED;
constant TAU_TAU_DIFF_PHI_LUT_SFIXED : calo_calo_diff_phi_lut_sfixed_array := CALO_CALO_DIFF_PHI_LUT_SFIXED;
constant TAU_PT_LUT_SFIXED : eg_pt_lut_sfixed_array := EG_PT_LUT_SFIXED;
constant EG_EG_COSH_DETA_LUT_SFIXED : calo_calo_cosh_deta_lut_sfixed_array := CALO_CALO_COSH_DETA_LUT_SFIXED;
constant EG_TAU_COSH_DETA_LUT_SFIXED : calo_calo_cosh_deta_lut_sfixed_array := CALO_CALO_COSH_DETA_LUT_SFIXED;
constant EG_JET_COSH_DETA_LUT_SFIXED : calo_calo_cosh_deta_lut_sfixed_array := CALO_CALO_COSH_DETA_LUT_SFIXED;
constant JET_EG_COSH_DETA_LUT_SFIXED : calo_calo_cosh_deta_lut_sfixed_array := CALO_CALO_COSH_DETA_LUT_SFIXED;
constant JET_JET_COSH_DETA_LUT_SFIXED : calo_calo_cosh_deta_lut_sfixed_array := CALO_CALO_COSH_DETA_LUT_SFIXED;
constant JET_TAU_COSH_DETA_LUT_SFIXED : calo_calo_cosh_deta_lut_sfixed_array := CALO_CALO_COSH_DETA_LUT_SFIXED;
constant TAU_EG_COSH_DETA_LUT_SFIXED : calo_calo_cosh_deta_lut_sfixed_array := CALO_CALO_COSH_DETA_LUT_SFIXED;
constant TAU_JET_COSH_DETA_LUT_SFIXED : calo_calo_cosh_deta_lut_sfixed_array := CALO_CALO_COSH_DETA_LUT_SFIXED;
constant TAU_TAU_COSH_DETA_LUT_SFIXED : calo_calo_cosh_deta_lut_sfixed_array := CALO_CALO_COSH_DETA_LUT_SFIXED;
constant EG_EG_COS_DPHI_LUT_SFIXED : calo_calo_cos_dphi_lut_sfixed_array := CALO_CALO_COS_DPHI_LUT_SFIXED;
constant EG_TAU_COS_DPHI_LUT_SFIXED : calo_calo_cos_dphi_lut_sfixed_array := CALO_CALO_COS_DPHI_LUT_SFIXED;
constant EG_JET_COS_DPHI_LUT_SFIXED : calo_calo_cos_dphi_lut_sfixed_array := CALO_CALO_COS_DPHI_LUT_SFIXED;
constant JET_EG_COS_DPHI_LUT_SFIXED : calo_calo_cos_dphi_lut_sfixed_array := CALO_CALO_COS_DPHI_LUT_SFIXED;
constant JET_JET_COS_DPHI_LUT_SFIXED : calo_calo_cos_dphi_lut_sfixed_array := CALO_CALO_COS_DPHI_LUT_SFIXED;
constant JET_TAU_COS_DPHI_LUT_SFIXED : calo_calo_cos_dphi_lut_sfixed_array := CALO_CALO_COS_DPHI_LUT_SFIXED;
constant TAU_EG_COS_DPHI_LUT_SFIXED : calo_calo_cos_dphi_lut_sfixed_array := CALO_CALO_COS_DPHI_LUT_SFIXED;
constant TAU_JET_COS_DPHI_LUT_SFIXED : calo_calo_cos_dphi_lut_sfixed_array := CALO_CALO_COS_DPHI_LUT_SFIXED;
constant TAU_TAU_COS_DPHI_LUT_SFIXED : calo_calo_cos_dphi_lut_sfixed_array := CALO_CALO_COS_DPHI_LUT_SFIXED;

end package;

