constant EG_EG_DIFF_ETA_LUT_SFIXED : calo_calo_diff_eta_lut_sfixed_array := CALO_CALO_DIFF_ETA_LUT_SFIXED;
constant EG_TAU_DIFF_ETA_LUT_SFIXED : calo_calo_diff_eta_lut_sfixed_array := CALO_CALO_DIFF_ETA_LUT_SFIXED;
constant EG_JET_DIFF_ETA_LUT_SFIXED : calo_calo_diff_eta_lut_sfixed_array := CALO_CALO_DIFF_ETA_LUT_SFIXED;
constant JET_EG_DIFF_ETA_LUT_SFIXED : calo_calo_diff_eta_lut_sfixed_array := CALO_CALO_DIFF_ETA_LUT_SFIXED;
constant JET_JET_DIFF_ETA_LUT_SFIXED : calo_calo_diff_eta_lut_sfixed_array := CALO_CALO_DIFF_ETA_LUT_SFIXED;
constant JET_TAU_DIFF_ETA_LUT_SFIXED : calo_calo_diff_eta_lut_sfixed_array := CALO_CALO_DIFF_ETA_LUT_SFIXED;
constant TAU_EG_DIFF_ETA_LUT_SFIXED : calo_calo_diff_eta_lut_sfixed_array := CALO_CALO_DIFF_ETA_LUT_SFIXED;
constant TAU_JET_DIFF_ETA_LUT_SFIXED : calo_calo_diff_eta_lut_sfixed_array := CALO_CALO_DIFF_ETA_LUT_SFIXED;
constant TAU_TAU_DIFF_ETA_LUT_SFIXED : calo_calo_diff_eta_lut_sfixed_array := CALO_CALO_DIFF_ETA_LUT_SFIXED;
constant EG_EG_DIFF_PHI_LUT_SFIXED : calo_calo_diff_phi_lut_sfixed_array := CALO_CALO_DIFF_PHI_LUT_SFIXED;
constant EG_TAU_DIFF_PHI_LUT_SFIXED : calo_calo_diff_phi_lut_sfixed_array := CALO_CALO_DIFF_PHI_LUT_SFIXED;
constant EG_JET_DIFF_PHI_LUT_SFIXED : calo_calo_diff_phi_lut_sfixed_array := CALO_CALO_DIFF_PHI_LUT_SFIXED;
constant JET_EG_DIFF_PHI_LUT_SFIXED : calo_calo_diff_phi_lut_sfixed_array := CALO_CALO_DIFF_PHI_LUT_SFIXED;
constant JET_JET_DIFF_PHI_LUT_SFIXED : calo_calo_diff_phi_lut_sfixed_array := CALO_CALO_DIFF_PHI_LUT_SFIXED;
constant JET_TAU_DIFF_PHI_LUT_SFIXED : calo_calo_diff_phi_lut_sfixed_array := CALO_CALO_DIFF_PHI_LUT_SFIXED;
constant TAU_EG_DIFF_PHI_LUT_SFIXED : calo_calo_diff_phi_lut_sfixed_array := CALO_CALO_DIFF_PHI_LUT_SFIXED;
constant TAU_JET_DIFF_PHI_LUT_SFIXED : calo_calo_diff_phi_lut_sfixed_array := CALO_CALO_DIFF_PHI_LUT_SFIXED;
constant TAU_TAU_DIFF_PHI_LUT_SFIXED : calo_calo_diff_phi_lut_sfixed_array := CALO_CALO_DIFF_PHI_LUT_SFIXED;
constant TAU_PT_LUT_SFIXED : eg_pt_lut_sfixed_array := EG_PT_LUT_SFIXED;
constant EG_EG_COSH_DETA_LUT_SFIXED : calo_calo_cosh_deta_lut_sfixed_array := CALO_CALO_COSH_DETA_LUT_SFIXED;
constant EG_TAU_COSH_DETA_LUT_SFIXED : calo_calo_cosh_deta_lut_sfixed_array := CALO_CALO_COSH_DETA_LUT_SFIXED;
constant EG_JET_COSH_DETA_LUT_SFIXED : calo_calo_cosh_deta_lut_sfixed_array := CALO_CALO_COSH_DETA_LUT_SFIXED;
constant JET_EG_COSH_DETA_LUT_SFIXED : calo_calo_cosh_deta_lut_sfixed_array := CALO_CALO_COSH_DETA_LUT_SFIXED;
constant JET_JET_COSH_DETA_LUT_SFIXED : calo_calo_cosh_deta_lut_sfixed_array := CALO_CALO_COSH_DETA_LUT_SFIXED;
constant JET_TAU_COSH_DETA_LUT_SFIXED : calo_calo_cosh_deta_lut_sfixed_array := CALO_CALO_COSH_DETA_LUT_SFIXED;
constant TAU_EG_COSH_DETA_LUT_SFIXED : calo_calo_cosh_deta_lut_sfixed_array := CALO_CALO_COSH_DETA_LUT_SFIXED;
constant TAU_JET_COSH_DETA_LUT_SFIXED : calo_calo_cosh_deta_lut_sfixed_array := CALO_CALO_COSH_DETA_LUT_SFIXED;
constant TAU_TAU_COSH_DETA_LUT_SFIXED : calo_calo_cosh_deta_lut_sfixed_array := CALO_CALO_COSH_DETA_LUT_SFIXED;
constant EG_EG_COS_DPHI_LUT_SFIXED : calo_calo_cos_dphi_lut_sfixed_array := CALO_CALO_COS_DPHI_LUT_SFIXED;
constant EG_TAU_COS_DPHI_LUT_SFIXED : calo_calo_cos_dphi_lut_sfixed_array := CALO_CALO_COS_DPHI_LUT_SFIXED;
constant EG_JET_COS_DPHI_LUT_SFIXED : calo_calo_cos_dphi_lut_sfixed_array := CALO_CALO_COS_DPHI_LUT_SFIXED;
constant JET_EG_COS_DPHI_LUT_SFIXED : calo_calo_cos_dphi_lut_sfixed_array := CALO_CALO_COS_DPHI_LUT_SFIXED;
constant JET_JET_COS_DPHI_LUT_SFIXED : calo_calo_cos_dphi_lut_sfixed_array := CALO_CALO_COS_DPHI_LUT_SFIXED;
constant JET_TAU_COS_DPHI_LUT_SFIXED : calo_calo_cos_dphi_lut_sfixed_array := CALO_CALO_COS_DPHI_LUT_SFIXED;
constant TAU_EG_COS_DPHI_LUT_SFIXED : calo_calo_cos_dphi_lut_sfixed_array := CALO_CALO_COS_DPHI_LUT_SFIXED;
constant TAU_JET_COS_DPHI_LUT_SFIXED : calo_calo_cos_dphi_lut_sfixed_array := CALO_CALO_COS_DPHI_LUT_SFIXED;
constant TAU_TAU_COS_DPHI_LUT_SFIXED : calo_calo_cos_dphi_lut_sfixed_array := CALO_CALO_COS_DPHI_LUT_SFIXED;

end package;

