library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all; -- for function "CONV_INTEGER"

use work.gtl_pkg.all;

package muon_phi_correction_pkg is

-- HB 2016-08-17: LUT was generated center values of pt and the formular: 2.677/pt**1.014 (pt [GeV] center value of bin). LUT values in bins.
type phi_correction_lut_array is array (0 to 2**(D_S_I_MUON.pt_high-D_S_I_MUON.pt_low)-1) of natural range 0 to 425;
constant PHI_CORRECTION_LUT : phi_correction_lut_array := (
0,	425,	329,	196,	139,	108,	88,	74,	64,	57,	51,	46,	42,	38,	35,	33,
31,	29,	27,	26,	24,	23,	22,	21,	20,	19,	19,	18,	17,	17,	16,	15,
15,	15,	14,	14,	13,	13,	13,	12,	12,	12,	11,	11,	11,	11,	10,	10,
10,	10,	9,	9,	9,	9,	9,	9,	8,	8,	8,	8,	8,	8,	8,	7,
7,	7,	7,	7,	7,	7,	7,	7,	7,	6,	6,	6,	6,	6,	6,	6,
6,	6,	6,	6,	6,	6,	5,	5,	5,	5,	5,	5,	5,	5,	5,	5,
5,	5,	5,	5,	5,	5,	5,	5,	4,	4,	4,	4,	4,	4,	4,	4,
4,	4,	4,	4,	4,	4,	4,	4,	4,	4,	4,	4,	4,	4,	4,	4,
4,	4,	4,	4,	4,	3,	3,	3,	3,	3,	3,	3,	3,	3,	3,	3,
3,	3,	3,	3,	3,	3,	3,	3,	3,	3,	3,	3,	3,	3,	3,	3,
3,	3,	3,	3,	3,	3,	3,	3,	3,	3,	3,	3,	3,	3,	3,	3,
3,	3,	3,	3,	3,	3,	3,	3,	3,	2,	2,	2,	2,	2,	2,	2,
2,	2,	2,	2,	2,	2,	2,	2,	2,	2,	2,	2,	2,	2,	2,	2,
2,	2,	2,	2,	2,	2,	2,	2,	2,	2,	2,	2,	2,	2,	2,	2,
2,	2,	2,	2,	2,	2,	2,	2,	2,	2,	2,	2,	2,	2,	2,	2,
2,	2,	2,	2,	2,	2,	2,	2,	2,	2,	2,	2,	2,	2,	2,	2,
2,	2,	2,	2,	2,	2,	2,	2,	2,	2,	2,	2,	2,	2,	2,	2,
2,	2,	2,	2,	2,	2,	2,	2,	2,	2,	2,	2,	2,	2,	2,	2,
2,	2,	2,	2,	2,	2,	2,	2,	2,	2,	2,	2,	2,	2,	2,	2,
2,	2,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,
1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,
1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,
1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,
1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,
1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,
1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,
1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,
1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,
1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,
1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,
1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,
1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1,	1
);

end package;
