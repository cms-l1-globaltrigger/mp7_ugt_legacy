library ieee;
use ieee.std_logic_1164.all;
package adt_test_sim_pkg is
constant ADT_ALGO_BIT: integer := 1;
constant ERROR_FILE_LOC: string := "/home/bergauer/github/cms-l1-globaltrigger/mp7_ugt_legacy/firmware/sim/adt_test/l1menu_adt_v6/module_2/error_file_L1_ADT_4000.txt";
end package;
