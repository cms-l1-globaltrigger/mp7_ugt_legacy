library ieee;
use ieee.std_logic_1164.all;
package adt_test_sim_pkg is
constant ADT_ALGO_BIT: integer := {{ALGO_BIT}};
constant ERROR_FILE_LOC: string := "{{ERR_FILE_LOC}}";
end package;
