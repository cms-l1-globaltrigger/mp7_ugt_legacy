-- Description:
-- Package for LUTS with sfixed format values.

-- Version history:
-- HB 2020-03-14: first design

library ieee;
use ieee.std_logic_1164.all;
-- use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
-- use ieee.numeric_std.all;
use ieee.fixed_pkg.all;

-- use work.lhc_data_pkg.all;
-- use work.math_pkg.all;
use work.gtl_pkg.all;

package sfixed_luts_pkg is

type calo_calo_diff_eta_lut_sfixed_array is array (0 to 2**MAX_CALO_ETA_BITS-1) of sfixed(5 downto -19);

constant CALO_CALO_DIFF_ETA_LUT_SFIXED : calo_calo_diff_eta_lut_sfixed_array := (
000000000000000000000000,
000000000101101000011100,
000000001011001000101101,
000000010000110001001001,
000000010110010001011010,
000000011011110001101010,
000000100001011010000111,
000000100111000010100011,
000000101100100010110100,
000000110010000011000100,
000000110111101011100001,
000000111101010011111101,
000001000010110100001110,
000001001000011100101011,
000001001101111100111011,
000001010011100101011000,
000001011001000101101000,
000001011110100101111000,
000001100100001110010101,
000001101001101110100101,
000001101111010111000010,
000001110100111111011111,
000001111010011111101111,
000010000000001000001100,
000010000101101000011100,
000010001011010000111001,
000010010000110001001001,
000010010110010001011010,
000010011011111001110110,
000010100001011010000111,
000010100111000010100011,
000010101100100010110100,
000010110010001011010000,
000010110111110011101101,
000010111101010011111101,
000011000010111100011010,
000011001000011100101011,
000011001110000101000111,
000011010011100101011000,
000011011001001101110100,
000011011110101110000101,
000011100100001110010101,
000011101001110110110010,
000011101111010111000010,
000011110100111111011111,
000011111010011111101111,
000100000000001000001100,
000100000101101000011100,
000100001011010000111001,
000100010000111001010110,
000100010110011001100110,
000100011011111001110110,
000100100001100010010011,
000100100111001010110000,
000100101100101011000000,
000100110010001011010000,
000100110111110011101101,
000100111101011100001010,
000101000010111100011010,
000101001000100100110111,
000101001110000101000111,
000101010011100101011000,
000101011001001101110100,
000101011110110110010001,
000101100100010110100001,
000101101001110110110010,
000101101111011111001110,
000101110101000111101011,
000101111010100111111011,
000110000000001000001100,
000110000101110000101000,
000110001011011001000101,
000110010000111001010110,
000110010110100001110010,
000110011100000010000011,
000110100001100010010011,
000110100111001010110000,
000110101100110011001100,
000110110010010011011101,
000110110111110011101101,
000110111101011100001010,
000111000011000100100110,
000111001000100100110111,
000111001110000101000111,
000111010011101101100100,
000111011001010110000001,
000111011110110110010001,
000111100100010110100001,
000111101001111110111110,
000111101111011111001110,
000111110101000111101011,
000111111010110000001000,
001000000000010000011000,
001000000101110000101000,
001000001011011001000101,
001000010000111001010110,
001000010110100001110010,
001000011100001010001111,
001000100001101010011111,
001000100111010010111100,
001000101100110011001100,
001000110010010011011101,
001000110111111011111001,
001000111101011100001010,
001001000011000100100110,
001001001000101101000011,
001001001110001101010011,
001001010011110101110000,
001001011001010110000001,
001001011110110110010001,
001001100100011110101110,
001001101010000111001010,
001001101111100111011011,
001001110101001111110111,
001001111010110000001000,
001010000000010000011000,
001010000101111000110101,
001010001011011001000101,
001010010001000001100010,
001010010110101001111110,
001010011100001010001111,
001010100001110010101100,
001010100111010010111100,
001010101100110011001100,
001010110010011011101001,
001010111000000100000110,
001010111101100100010110,
001011000011001100110011,
001011001000101101000011,
001011001110001101010011,
001011010011110101110000,
001011011001010110000001,
001011011110111110011101,
001011100100100110111010,
001011101010000111001010,
001011101111101111100111,
001011110101001111110111,
001011111010110000001000,
001100000000011000100100,
001100000110000001000001,
001100001011100001010001,
001100010001001001101110,
001100010110101001111110,
001100011100001010001111,
001100100001110010101100,
001100100111010010111100,
001100101100111011011001,
001100110010100011110101,
001100111000000100000110,
001100111101101100100010,
001101000011001100110011,
001101001000101101000011,
001101001110010101100000,
001101010011111101111100,
001101011001011110001101,
001101011111000110101001,
001101100100100110111010,
001101101010000111001010,
001101101111101111100111,
001101110101001111110111,
001101111010111000010100,
001110000000100000110001,
001110000110000001000001,
001110001011101001011110,
001110010001001001101110,
001110010110101001111110,
001110011100010010011011,
001110100001110010101100,
001110100111011011001000,
001110101101000011100101,
001110110010100011110101,
001110111000000100000110,
001110111101101100100010,
001111000011001100110011,
001111001000110101001111,
001111001110011101101100,
001111010011111101111100,
001111011001100110011001,
001111011111000110101001,
001111100100100110111010,
001111101010001111010111,
001111101111101111100111,
001111110101011000000100,
001111111011000000100000,
010000000000100000110001,
010000000110000001000001,
010000001011101001011110,
010000010001001001101110,
010000010110110010001011,
010000011100010010011011,
010000100001111010111000,
010000100111011011001000,
010000101101000011100101,
010000110010101100000010,
010000111000001100010010,
010000111101110100101111,
010001000011010100111111,
010001001000111101011100,
010001001110011101101100,
010001010100000110001001,
010001011001100110011001,
010001011111001110110110,
010001100100101111000110,
010001101010001111010111,
010001101111110111110011,
010001110101011000000100,
010001111011000000100000,
010010000000101000111101,
010010000110001001001101,
010010001011110001101010,
010010010001010001111010,
010010010110111010010111,
010010011100011010100111,
010010100010000011000100,
010010100111100011010100,
010010101101001011110001,
010010110010101100000010,
010010111000001100010010,
010010111101110100101111,
010011000011010100111111,
010011001000111101011100,
010011001110100101111000,
010011010100000110001001,
010011011001101110100101,
010011011111001110110110,
010011100100110111010010,
010011101010010111100011,
010011101111111111111111,
010011110101100000010000,
010011111011001000101101,
000000000000000000000000,
000000000000000000000000,
000000000000000000000000,
000000000000000000000000,
000000000000000000000000,
000000000000000000000000,
000000000000000000000000,
000000000000000000000000,
000000000000000000000000,
000000000000000000000000,
000000000000000000000000,
000000000000000000000000,
000000000000000000000000,
000000000000000000000000,
000000000000000000000000,
000000000000000000000000,
000000000000000000000000,
000000000000000000000000,
000000000000000000000000,
000000000000000000000000,
000000000000000000000000,
000000000000000000000000,
000000000000000000000000,
000000000000000000000000,
000000000000000000000000,
000000000000000000000000
);

constant EG_EG_DIFF_ETA_LUT_SFIXED : calo_calo_diff_eta_lut_array := CALO_CALO_DIFF_ETA_LUT_SFIXED;
constant EG_TAU_DIFF_ETA_LUT_SFIXED : calo_calo_diff_eta_lut_array := CALO_CALO_DIFF_ETA_LUT_SFIXED;
constant EG_JET_DIFF_ETA_LUT_SFIXED : calo_calo_diff_eta_lut_array := CALO_CALO_DIFF_ETA_LUT_SFIXED;
constant JET_EG_DIFF_ETA_LUT_SFIXED : calo_calo_diff_eta_lut_array := CALO_CALO_DIFF_ETA_LUT_SFIXED;
constant JET_JET_DIFF_ETA_LUT_SFIXED : calo_calo_diff_eta_lut_array := CALO_CALO_DIFF_ETA_LUT_SFIXED;
constant JET_TAU_DIFF_ETA_LUT_SFIXED : calo_calo_diff_eta_lut_array := CALO_CALO_DIFF_ETA_LUT_SFIXED;
constant TAU_EG_DIFF_ETA_LUT_SFIXED : calo_calo_diff_eta_lut_array := CALO_CALO_DIFF_ETA_LUT_SFIXED;
constant TAU_JET_DIFF_ETA_LUT_SFIXED : calo_calo_diff_eta_lut_array := CALO_CALO_DIFF_ETA_LUT_SFIXED;
constant TAU_TAU_DIFF_ETA_LUT_SFIXED : calo_calo_diff_eta_lut_array := CALO_CALO_DIFF_ETA_LUT_SFIXED;

type calo_calo_diff_phi_lut_sfixed_array is array (0 to 2**MAX_CALO_PHI_BITS-1) of sfixed(4 downto -19);

constant CALO_CALO_DIFF_PHI_LUT_SFIXED : calo_calo_diff_phi_lut_sfixed_array := (
00000000000000000000000,
00000000101101000011100,
00000001011001000101101,
00000010000110001001001,
00000010110011001100110,
00000011011111001110110,
00000100001100010010011,
00000100111000010100011,
00000101100101011000000,
00000110010010011011101,
00000110111110011101101,
00000111101011100001010,
00001000011000100100110,
00001001000100100110111,
00001001110001101010011,
00001010011101101100100,
00001011001010110000001,
00001011110111110011101,
00001100100011110101110,
00001101010000111001010,
00001101111101111100111,
00001110101001111110111,
00001111010111000010100,
00010000000100000110001,
00010000110000001000001,
00010001011101001011110,
00010010001001001101110,
00010010110110010001011,
00010011100011010100111,
00010100001111010111000,
00010100111100011010100,
00010101101001011110001,
00010110010101100000010,
00010111000010100011110,
00010111101111100111011,
00011000011011101001011,
00011001001000101101000,
00011001110100101111000,
00011010100001110010101,
00011011001110110110010,
00011011111010111000010,
00011100100111111011111,
00011101010100111111011,
00011110000001000001100,
00011110101110000101000,
00011111011010000111001,
00100000000111001010110,
00100000110100001110010,
00100001100000010000011,
00100010001101010011111,
00100010111010010111100,
00100011100110011001100,
00100100010011011101001,
00100101000000100000110,
00100101101100100010110,
00100110011001100110011,
00100111000101101000011,
00100111110010101100000,
00101000011111101111100,
00101001001011110001101,
00101001111000110101001,
00101010100101111000110,
00101011010001111010111,
00101011111110111110011,
00101100101100000010000,
00101101011000000100000,
00101110000101000111101,
00101110110001001001101,
00101111011110001101010,
00110000001011010000111,
00110000110111010010111,
00110001100100010110100,
00110010010001011010000,
00110010111101011100001,
00110011101010011111101,
00110100010110100001110,
00110101000011100101011,
00110101110000101000111,
00110110011100101011000,
00110111001001101110100,
00110111110110110010001,
00111000100010110100001,
00111001001111110111110,
00111001111100111011011,
00111010101000111101011,
00111011010110000001000,
00111100000010000011000,
00111100101111000110101,
00111101011100001010001,
00111110001000001100010,
00111110110101001111110,
00111111100010010011011,
01000000001110010101100,
01000000111011011001000,
01000001101000011100101,
01000010010100011110101,
01000011000001100010010,
01000011101101100100010,
01000100011010100111111,
01000101000111101011100,
01000101110011101101100,
01000110100000110001001,
01000111001101110100101,
01000111111001110110110,
01001000100110111010010,
01001001010010111100011,
01001001111111111111111,
01001010101101000011100,
01001011011001000101101,
01001100000110001001001,
01001100110011001100110,
01001101011111001110110,
01001110001100010010011,
01001110111001010110000,
01001111100101011000000,
01010000010010011011101,
01010000111110011101101,
01010001101011100001010,
01010010011000100100110,
01010011000100100110111,
01010011110001101010011,
01010100011110101110000,
01010101001010110000001,
01010101110111110011101,
01010110100100110111010,
01010111010000111001010,
01010111111101111100111,
01011000101001111110111,
01011001010111000010100,
01011010000100000110001,
01011010110000001000001,
01011011011101001011110,
01011100001010001111010,
01011100110110010001011,
01011101100011010100111,
01011110001111010111000,
01011110111100011010100,
01011111101001011110001,
01100000010101100000010,
01100001000010100011110,
01100001101111100111011,
01100010011011101001011,
01100011001000101101000,
01100011110101110000101,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000
);

constant EG_EG_DIFF_PHI_LUT_SFIXED : calo_calo_diff_phi_lut_array := CALO_CALO_DIFF_PHI_LUT_SFIXED;
constant EG_TAU_DIFF_PHI_LUT_SFIXED : calo_calo_diff_phi_lut_array := CALO_CALO_DIFF_PHI_LUT_SFIXED;
constant EG_JET_DIFF_PHI_LUT_SFIXED : calo_calo_diff_phi_lut_array := CALO_CALO_DIFF_PHI_LUT_SFIXED;
constant JET_EG_DIFF_PHI_LUT_SFIXED : calo_calo_diff_phi_lut_array := CALO_CALO_DIFF_PHI_LUT_SFIXED;
constant JET_JET_DIFF_PHI_LUT_SFIXED : calo_calo_diff_phi_lut_array := CALO_CALO_DIFF_PHI_LUT_SFIXED;
constant JET_TAU_DIFF_PHI_LUT_SFIXED : calo_calo_diff_phi_lut_array := CALO_CALO_DIFF_PHI_LUT_SFIXED;
constant TAU_EG_DIFF_PHI_LUT_SFIXED : calo_calo_diff_phi_lut_array := CALO_CALO_DIFF_PHI_LUT_SFIXED;
constant TAU_JET_DIFF_PHI_LUT_SFIXED : calo_calo_diff_phi_lut_array := CALO_CALO_DIFF_PHI_LUT_SFIXED;
constant TAU_TAU_DIFF_PHI_LUT_SFIXED : calo_calo_diff_phi_lut_array := CALO_CALO_DIFF_PHI_LUT_SFIXED;

-- muon-muon differences LUTs
type muon_muon_diff_eta_lut_array is array (0 to 2**(MUON_ETA_HIGH-MUON_ETA_LOW+1)-1) of sfixed(4 downto -19);

constant MU_MU_DIFF_ETA_LUT_SFIXED : muon_muon_diff_eta_lut_array := (
00000000000000000000000,
00000000001011010000111,
00000000010110100001110,
00000000100001110010101,
00000000101101000011100,
00000000110111010010111,
00000001000010100011110,
00000001001101110100101,
00000001011001000101101,
00000001100100010110100,
00000001101111100111011,
00000001111010111000010,
00000010000110001001001,
00000010010000011000100,
00000010011011101001011,
00000010100110111010010,
00000010110010001011010,
00000010111101011100001,
00000011001000101101000,
00000011010011111101111,
00000011011110001101010,
00000011101001011110001,
00000011110100101111000,
00000011111111111111111,
00000100001011010000111,
00000100010110100001110,
00000100100001110010101,
00000100101101000011100,
00000100111000010100011,
00000101000010100011110,
00000101001101110100101,
00000101011001000101101,
00000101100100010110100,
00000101101111100111011,
00000101111010111000010,
00000110000110001001001,
00000110010000011000100,
00000110011011101001011,
00000110100110111010010,
00000110110010001011010,
00000110111101011100001,
00000111001000101101000,
00000111010011111101111,
00000111011111001110110,
00000111101010011111101,
00000111110100101111000,
00000111111111111111111,
00001000001011010000111,
00001000010110100001110,
00001000100001110010101,
00001000101101000011100,
00001000111000010100011,
00001001000011100101011,
00001001001101110100101,
00001001011001000101101,
00001001100100010110100,
00001001101111100111011,
00001001111010111000010,
00001010000110001001001,
00001010010001011010000,
00001010011100101011000,
00001010100110111010010,
00001010110010001011010,
00001010111101011100001,
00001011001000101101000,
00001011010011111101111,
00001011011111001110110,
00001011101010011111101,
00001011110100101111000,
00001011111111111111111,
00001100001011010000111,
00001100010110100001110,
00001100100001110010101,
00001100101101000011100,
00001100111000010100011,
00001101000011100101011,
00001101001101110100101,
00001101011001000101101,
00001101100100010110100,
00001101101111100111011,
00001101111010111000010,
00001110000110001001001,
00001110010001011010000,
00001110011100101011000,
00001110100111111011111,
00001110110010001011010,
00001110111101011100001,
00001111001000101101000,
00001111010011111101111,
00001111011111001110110,
00001111101010011111101,
00001111110101110000101,
00010000000001000001100,
00010000001011010000111,
00010000010110100001110,
00010000100001110010101,
00010000101101000011100,
00010000111000010100011,
00010001000011100101011,
00010001001110110110010,
00010001011010000111001,
00010001100100010110100,
00010001101111100111011,
00010001111010111000010,
00010010000110001001001,
00010010010001011010000,
00010010011100101011000,
00010010100111111011111,
00010010110010001011010,
00010010111101011100001,
00010011001000101101000,
00010011010011111101111,
00010011011111001110110,
00010011101010011111101,
00010011110101110000101,
00010100000001000001100,
00010100001011010000111,
00010100010110100001110,
00010100100001110010101,
00010100101101000011100,
00010100111000010100011,
00010101000011100101011,
00010101001110110110010,
00010101011010000111001,
00010101100100010110100,
00010101101111100111011,
00010101111010111000010,
00010110000110001001001,
00010110010001011010000,
00010110011100101011000,
00010110100111111011111,
00010110110011001100110,
00010110111110011101101,
00010111001000101101000,
00010111010011111101111,
00010111011111001110110,
00010111101010011111101,
00010111110101110000101,
00011000000001000001100,
00011000001100010010011,
00011000010111100011010,
00011000100001110010101,
00011000101101000011100,
00011000111000010100011,
00011001000011100101011,
00011001001110110110010,
00011001011010000111001,
00011001100101011000000,
00011001110000101000111,
00011001111010111000010,
00011010000110001001001,
00011010010001011010000,
00011010011100101011000,
00011010100111111011111,
00011010110011001100110,
00011010111110011101101,
00011011001001101110100,
00011011010011111101111,
00011011011111001110110,
00011011101010011111101,
00011011110101110000101,
00011100000001000001100,
00011100001100010010011,
00011100010111100011010,
00011100100001110010101,
00011100101101000011100,
00011100111000010100011,
00011101000011100101011,
00011101001110110110010,
00011101011010000111001,
00011101100101011000000,
00011101110000101000111,
00011101111010111000010,
00011110000110001001001,
00011110010001011010000,
00011110011100101011000,
00011110100111111011111,
00011110110011001100110,
00011110111110011101101,
00011111001001101110100,
00011111010011111101111,
00011111011111001110110,
00011111101010011111101,
00011111110101110000101,
00100000000001000001100,
00100000001100010010011,
00100000010111100011010,
00100000100010110100001,
00100000101101000011100,
00100000111000010100011,
00100001000011100101011,
00100001001110110110010,
00100001011010000111001,
00100001100101011000000,
00100001110000101000111,
00100001111011111001110,
00100010000111001010110,
00100010010001011010000,
00100010011100101011000,
00100010100111111011111,
00100010110011001100110,
00100010111110011101101,
00100011001001101110100,
00100011010100111111011,
00100011011111001110110,
00100011101010011111101,
00100011110101110000101,
00100100000001000001100,
00100100001100010010011,
00100100010111100011010,
00100100100010110100001,
00100100101110000101000,
00100100111001010110000,
00100101000011100101011,
00100101001110110110010,
00100101011010000111001,
00100101100101011000000,
00100101110000101000111,
00100101111011111001110,
00100110000111001010110,
00100110010001011010000,
00100110011100101011000,
00100110100111111011111,
00100110110011001100110,
00100110111110011101101,
00100111001001101110100,
00100111010100111111011,
00100111100000010000011,
00100111101011100001010,
00100111110101110000101,
00101000000001000001100,
00101000001100010010011,
00101000010111100011010,
00101000100010110100001,
00101000101110000101000,
00101000111001010110000,
00101001000100100110111,
00101001001110110110010,
00101001011010000111001,
00101001100101011000000,
00101001110000101000111,
00101001111011111001110,
00101010000111001010110,
00101010010010011011101,
00101010011100101011000,
00101010100111111011111,
00101010110011001100110,
00101010111110011101101,
00101011001001101110100,
00101011010100111111011,
00101011100000010000011,
00101011101011100001010,
00101011110110110010001,
00101100000001000001100,
00101100001100010010011,
00101100010111100011010,
00101100100010110100001,
00101100101110000101000,
00101100111001010110000,
00101101000100100110111,
00101101001110110110010,
00101101011010000111001,
00101101100101011000000,
00101101110000101000111,
00101101111011111001110,
00101110000111001010110,
00101110010010011011101,
00101110011101101100100,
00101110101000111101011,
00101110110011001100110,
00101110111110011101101,
00101111001001101110100,
00101111010100111111011,
00101111100000010000011,
00101111101011100001010,
00101111110110110010001,
00110000000001000001100,
00110000001100010010011,
00110000010111100011010,
00110000100010110100001,
00110000101110000101000,
00110000111001010110000,
00110001000100100110111,
00110001001111110111110,
00110001011011001000101,
00110001100101011000000,
00110001110000101000111,
00110001111011111001110,
00110010000111001010110,
00110010010010011011101,
00110010011101101100100,
00110010101000111101011,
00110010110100001110010,
00110010111110011101101,
00110011001001101110100,
00110011010100111111011,
00110011100000010000011,
00110011101011100001010,
00110011110110110010001,
00110100000010000011000,
00110100001100010010011,
00110100010111100011010,
00110100100010110100001,
00110100101110000101000,
00110100111001010110000,
00110101000100100110111,
00110101001111110111110,
00110101011011001000101,
00110101100110011001100,
00110101110000101000111,
00110101111011111001110,
00110110000111001010110,
00110110010010011011101,
00110110011101101100100,
00110110101000111101011,
00110110110100001110010,
00110110111110011101101,
00110111001001101110100,
00110111010100111111011,
00110111100000010000011,
00110111101011100001010,
00110111110110110010001,
00111000000010000011000,
00111000001101010011111,
00111000011000100100110,
00111000100010110100001,
00111000101110000101000,
00111000111001010110000,
00111001000100100110111,
00111001001111110111110,
00111001011011001000101,
00111001100110011001100,
00111001110000101000111,
00111001111011111001110,
00111010000111001010110,
00111010010010011011101,
00111010011101101100100,
00111010101000111101011,
00111010110100001110010,
00111010111111011111001,
00111011001010110000001,
00111011010100111111011,
00111011100000010000011,
00111011101011100001010,
00111011110110110010001,
00111100000010000011000,
00111100001101010011111,
00111100011000100100110,
00111100100010110100001,
00111100101110000101000,
00111100111001010110000,
00111101000100100110111,
00111101001111110111110,
00111101011011001000101,
00111101100110011001100,
00111101110001101010011,
00111101111011111001110,
00111110000111001010110,
00111110010010011011101,
00111110011101101100100,
00111110101000111101011,
00111110110100001110010,
00111110111111011111001,
00111111001010110000001,
00111111010110000001000,
00111111100000010000011,
00111111101011100001010,
00111111110110110010001,
01000000000010000011000,
01000000001101010011111,
01000000011000100100110,
01000000100011110101110,
01000000101110000101000,
01000000111001010110000,
01000001000100100110111,
01000001001111110111110,
01000001011011001000101,
01000001100110011001100,
01000001110001101010011,
01000001111100111011011,
01000010000111001010110,
01000010010010011011101,
01000010011101101100100,
01000010101000111101011,
01000010110100001110010,
01000010111111011111001,
01000011001010110000001,
01000011010110000001000,
01000011100001010001111,
01000011101011100001010,
01000011110110110010001,
01000100000010000011000,
01000100001101010011111,
01000100011000100100110,
01000100100011110101110,
01000100101111000110101,
01000100111010010111100,
01000101000100100110111,
01000101001111110111110,
01000101011011001000101,
01000101100110011001100,
01000101110001101010011,
01000101111100111011011,
01000110001000001100010,
01000110010010011011101,
01000110011101101100100,
01000110101000111101011,
01000110110100001110010,
01000110111111011111001,
01000111001010110000001,
01000111010110000001000,
01000111100001010001111,
01000111101011100001010,
01000111110110110010001,
01001000000010000011000,
01001000001101010011111,
01001000011000100100110,
01001000100011110101110,
01001000101111000110101,
01001000111010010111100,
01001001000101101000011,
01001001001111110111110,
01001001011011001000101,
01001001100110011001100,
01001001110001101010011,
01001001111100111011011,
01001010001000001100010,
01001010010011011101001,
01001010011110101110000,
01001010101000111101011,
01001010110100001110010,
01001010111111011111001,
01001011001010110000001,
01001011010110000001000,
01001011100001010001111,
01001011101100100010110,
01001011110110110010001,
01001100000010000011000,
01001100001101010011111,
01001100011000100100110,
01001100100011110101110,
01001100101111000110101,
01001100111010010111100,
01001101000101101000011,
01001101010000111001010,
01001101011011001000101,
01001101100110011001100,
01001101110001101010011,
01001101111100111011011,
01001110001000001100010,
01001110010011011101001,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000
);

type muon_muon_diff_phi_lut_array is array (0 to 2**(MUON_PHI_HIGH-MUON_PHI_LOW+1)-1) of sfixed(4 downto -19);

constant MU_MU_DIFF_PHI_LUT_SFIXED : muon_muon_diff_phi_lut_array := (
00000000000000000000000,
00000000001011010000111,
00000000010110100001110,
00000000100001110010101,
00000000101101000011100,
00000000111000010100011,
00000001000010100011110,
00000001001101110100101,
00000001011001000101101,
00000001100100010110100,
00000001101111100111011,
00000001111010111000010,
00000010000110001001001,
00000010010001011010000,
00000010011100101011000,
00000010100111111011111,
00000010110011001100110,
00000010111101011100001,
00000011001000101101000,
00000011010011111101111,
00000011011111001110110,
00000011101010011111101,
00000011110101110000101,
00000100000001000001100,
00000100001100010010011,
00000100010111100011010,
00000100100010110100001,
00000100101110000101000,
00000100111000010100011,
00000101000011100101011,
00000101001110110110010,
00000101011010000111001,
00000101100101011000000,
00000101110000101000111,
00000101111011111001110,
00000110000111001010110,
00000110010010011011101,
00000110011101101100100,
00000110101000111101011,
00000110110011001100110,
00000110111110011101101,
00000111001001101110100,
00000111010100111111011,
00000111100000010000011,
00000111101011100001010,
00000111110110110010001,
00001000000010000011000,
00001000001101010011111,
00001000011000100100110,
00001000100011110101110,
00001000101110000101000,
00001000111001010110000,
00001001000100100110111,
00001001001111110111110,
00001001011011001000101,
00001001100110011001100,
00001001110001101010011,
00001001111100111011011,
00001010001000001100010,
00001010010011011101001,
00001010011101101100100,
00001010101000111101011,
00001010110100001110010,
00001010111111011111001,
00001011001010110000001,
00001011010110000001000,
00001011100001010001111,
00001011101100100010110,
00001011110111110011101,
00001100000011000100100,
00001100001110010101100,
00001100011000100100110,
00001100100011110101110,
00001100101111000110101,
00001100111010010111100,
00001101000101101000011,
00001101010000111001010,
00001101011100001010001,
00001101100111011011001,
00001101110010101100000,
00001101111101111100111,
00001110001001001101110,
00001110010011011101001,
00001110011110101110000,
00001110101001111110111,
00001110110101001111110,
00001111000000100000110,
00001111001011110001101,
00001111010111000010100,
00001111100010010011011,
00001111101101100100010,
00001111111000110101001,
00010000000100000110001,
00010000001110010101100,
00010000011001100110011,
00010000100100110111010,
00010000110000001000001,
00010000111011011001000,
00010001000110101001111,
00010001010001111010111,
00010001011101001011110,
00010001101000011100101,
00010001110011101101100,
00010001111110111110011,
00010010001001001101110,
00010010010100011110101,
00010010011111101111100,
00010010101011000000100,
00010010110110010001011,
00010011000001100010010,
00010011001100110011001,
00010011011000000100000,
00010011100011010100111,
00010011101110100101111,
00010011111001110110110,
00010100000100000110001,
00010100001111010111000,
00010100011010100111111,
00010100100101111000110,
00010100110001001001101,
00010100111100011010100,
00010101000111101011100,
00010101010010111100011,
00010101011110001101010,
00010101101001011110001,
00010101110100101111000,
00010101111110111110011,
00010110001010001111010,
00010110010101100000010,
00010110100000110001001,
00010110101100000010000,
00010110110111010010111,
00010111000010100011110,
00010111001101110100101,
00010111011001000101101,
00010111100100010110100,
00010111101111100111011,
00010111111001110110110,
00011000000101000111101,
00011000010000011000100,
00011000011011101001011,
00011000100110111010010,
00011000110010001011010,
00011000111101011100001,
00011001001000101101000,
00011001010011111101111,
00011001011111001110110,
00011001101010011111101,
00011001110100101111000,
00011001111111111111111,
00011010001011010000111,
00011010010110100001110,
00011010100001110010101,
00011010101101000011100,
00011010111000010100011,
00011011000011100101011,
00011011001110110110010,
00011011011010000111001,
00011011100101011000000,
00011011101111100111011,
00011011111010111000010,
00011100000110001001001,
00011100010001011010000,
00011100011100101011000,
00011100100111111011111,
00011100110011001100110,
00011100111110011101101,
00011101001001101110100,
00011101010100111111011,
00011101100000010000011,
00011101101010011111101,
00011101110101110000101,
00011110000001000001100,
00011110001100010010011,
00011110010111100011010,
00011110100010110100001,
00011110101110000101000,
00011110111001010110000,
00011111000100100110111,
00011111001111110111110,
00011111011010000111001,
00011111100101011000000,
00011111110000101000111,
00011111111011111001110,
00100000000111001010110,
00100000010010011011101,
00100000011101101100100,
00100000101000111101011,
00100000110100001110010,
00100000111111011111001,
00100001001010110000001,
00100001010100111111011,
00100001100000010000011,
00100001101011100001010,
00100001110110110010001,
00100010000010000011000,
00100010001101010011111,
00100010011000100100110,
00100010100011110101110,
00100010101111000110101,
00100010111010010111100,
00100011000101101000011,
00100011001111110111110,
00100011011011001000101,
00100011100110011001100,
00100011110001101010011,
00100011111100111011011,
00100100001000001100010,
00100100010011011101001,
00100100011110101110000,
00100100101001111110111,
00100100110101001111110,
00100101000000100000110,
00100101001010110000001,
00100101010110000001000,
00100101100001010001111,
00100101101100100010110,
00100101110111110011101,
00100110000011000100100,
00100110001110010101100,
00100110011001100110011,
00100110100100110111010,
00100110110000001000001,
00100110111011011001000,
00100111000101101000011,
00100111010000111001010,
00100111011100001010001,
00100111100111011011001,
00100111110010101100000,
00100111111101111100111,
00101000001001001101110,
00101000010100011110101,
00101000011111101111100,
00101000101011000000100,
00101000110110010001011,
00101001000000100000110,
00101001001011110001101,
00101001010111000010100,
00101001100010010011011,
00101001101101100100010,
00101001111000110101001,
00101010000100000110001,
00101010001111010111000,
00101010011010100111111,
00101010100101111000110,
00101010110001001001101,
00101010111011011001000,
00101011000110101001111,
00101011010001111010111,
00101011011101001011110,
00101011101000011100101,
00101011110011101101100,
00101011111110111110011,
00101100001010001111010,
00101100010101100000010,
00101100100000110001001,
00101100101100000010000,
00101100110110010001011,
00101101000001100010010,
00101101001100110011001,
00101101011000000100000,
00101101100011010100111,
00101101101110100101111,
00101101111001110110110,
00101110000101000111101,
00101110010000011000100,
00101110011011101001011,
00101110100110111010010,
00101110110001001001101,
00101110111100011010100,
00101111000111101011100,
00101111010010111100011,
00101111011110001101010,
00101111101001011110001,
00101111110100101111000,
00110000000000000000000,
00110000001011010000111,
00110000010110100001110,
00110000100001110010101,
00110000101100000010000,
00110000110111010010111,
00110001000010100011110,
00110001001101110100101,
00110001011001000101101,
00110001100100010110100,
00110001101111100111011,
00110001111010111000010,
00110010000110001001001,
00110010010001011010000,
00110010011100101011000,
00110010100110111010010,
00110010110010001011010,
00110010111101011100001,
00110011001000101101000,
00110011010011111101111,
00110011011111001110110,
00110011101010011111101,
00110011110101110000101,
00110100000001000001100,
00110100001100010010011,
00110100010110100001110,
00110100100001110010101,
00110100101101000011100,
00110100111000010100011,
00110101000011100101011,
00110101001110110110010,
00110101011010000111001,
00110101100101011000000,
00110101110000101000111,
00110101111011111001110,
00110110000111001010110,
00110110010001011010000,
00110110011100101011000,
00110110100111111011111,
00110110110011001100110,
00110110111110011101101,
00110111001001101110100,
00110111010100111111011,
00110111100000010000011,
00110111101011100001010,
00110111110110110010001,
00111000000010000011000,
00111000001100010010011,
00111000010111100011010,
00111000100010110100001,
00111000101110000101000,
00111000111001010110000,
00111001000100100110111,
00111001001111110111110,
00111001011011001000101,
00111001100110011001100,
00111001110001101010011,
00111001111100111011011,
00111010000111001010110,
00111010010010011011101,
00111010011101101100100,
00111010101000111101011,
00111010110100001110010,
00111010111111011111001,
00111011001010110000001,
00111011010110000001000,
00111011100001010001111,
00111011101100100010110,
00111011110111110011101,
00111100000010000011000,
00111100001101010011111,
00111100011000100100110,
00111100100011110101110,
00111100101111000110101,
00111100111010010111100,
00111101000101101000011,
00111101010000111001010,
00111101011100001010001,
00111101100111011011001,
00111101110010101100000,
00111101111100111011011,
00111110001000001100010,
00111110010011011101001,
00111110011110101110000,
00111110101001111110111,
00111110110101001111110,
00111111000000100000110,
00111111001011110001101,
00111111010111000010100,
00111111100010010011011,
00111111101101100100010,
00111111110111110011101,
01000000000011000100100,
01000000001110010101100,
01000000011001100110011,
01000000100100110111010,
01000000110000001000001,
01000000111011011001000,
01000001000110101001111,
01000001010001111010111,
01000001011101001011110,
01000001101000011100101,
01000001110010101100000,
01000001111101111100111,
01000010001001001101110,
01000010010100011110101,
01000010011111101111100,
01000010101011000000100,
01000010110110010001011,
01000011000001100010010,
01000011001100110011001,
01000011011000000100000,
01000011100011010100111,
01000011101101100100010,
01000011111000110101001,
01000100000100000110001,
01000100001111010111000,
01000100011010100111111,
01000100100101111000110,
01000100110001001001101,
01000100111100011010100,
01000101000111101011100,
01000101010010111100011,
01000101011110001101010,
01000101101000011100101,
01000101110011101101100,
01000101111110111110011,
01000110001010001111010,
01000110010101100000010,
01000110100000110001001,
01000110101100000010000,
01000110110111010010111,
01000111000010100011110,
01000111001101110100101,
01000111011000000100000,
01000111100011010100111,
01000111101110100101111,
01000111111001110110110,
01001000000101000111101,
01001000010000011000100,
01001000011011101001011,
01001000100110111010010,
01001000110010001011010,
01001000111101011100001,
01001001001000101101000,
01001001010010111100011,
01001001011110001101010,
01001001101001011110001,
01001001110100101111000,
01001001111111111111111,
01001010001011010000111,
01001010010110100001110,
01001010100001110010101,
01001010101101000011100,
01001010111000010100011,
01001011000011100101011,
01001011001101110100101,
01001011011001000101101,
01001011100100010110100,
01001011101111100111011,
01001011111010111000010,
01001100000110001001001,
01001100010001011010000,
01001100011100101011000,
01001100100111111011111,
01001100110011001100110,
01001100111110011101101,
01001101001000101101000,
01001101010011111101111,
01001101011111001110110,
01001101101010011111101,
01001101110101110000101,
01001110000001000001100,
01001110001100010010011,
01001110010111100011010,
01001110100010110100001,
01001110101110000101000,
01001110111001010110000,
01001111000011100101011,
01001111001110110110010,
01001111011010000111001,
01001111100101011000000,
01001111110000101000111,
01001111111011111001110,
01010000000111001010110,
01010000010010011011101,
01010000011101101100100,
01010000101000111101011,
01010000110100001110010,
01010000111110011101101,
01010001001001101110100,
01010001010100111111011,
01010001100000010000011,
01010001101011100001010,
01010001110110110010001,
01010010000010000011000,
01010010001101010011111,
01010010011000100100110,
01010010100011110101110,
01010010101111000110101,
01010010111001010110000,
01010011000100100110111,
01010011001111110111110,
01010011011011001000101,
01010011100110011001100,
01010011110001101010011,
01010011111100111011011,
01010100001000001100010,
01010100010011011101001,
01010100011110101110000,
01010100101001111110111,
01010100110100001110010,
01010100111111011111001,
01010101001010110000001,
01010101010110000001000,
01010101100001010001111,
01010101101100100010110,
01010101110111110011101,
01010110000011000100100,
01010110001110010101100,
01010110011001100110011,
01010110100100110111010,
01010110101111000110101,
01010110111010010111100,
01010111000101101000011,
01010111010000111001010,
01010111011100001010001,
01010111100111011011001,
01010111110010101100000,
01010111111101111100111,
01011000001001001101110,
01011000010100011110101,
01011000011111101111100,
01011000101001111110111,
01011000110101001111110,
01011001000000100000110,
01011001001011110001101,
01011001010111000010100,
01011001100010010011011,
01011001101101100100010,
01011001111000110101001,
01011010000100000110001,
01011010001111010111000,
01011010011010100111111,
01011010100100110111010,
01011010110000001000001,
01011010111011011001000,
01011011000110101001111,
01011011010001111010111,
01011011011101001011110,
01011011101000011100101,
01011011110011101101100,
01011011111110111110011,
01011100001010001111010,
01011100010100011110101,
01011100011111101111100,
01011100101011000000100,
01011100110110010001011,
01011101000001100010010,
01011101001100110011001,
01011101011000000100000,
01011101100011010100111,
01011101101110100101111,
01011101111001110110110,
01011110000101000111101,
01011110001111010111000,
01011110011010100111111,
01011110100101111000110,
01011110110001001001101,
01011110111100011010100,
01011111000111101011100,
01011111010010111100011,
01011111011110001101010,
01011111101001011110001,
01011111110100101111000,
01100000000000000000000,
01100000001010001111010,
01100000010101100000010,
01100000100000110001001,
01100000101100000010000,
01100000110111010010111,
01100001000010100011110,
01100001001101110100101,
01100001011001000101101,
01100001100100010110100,
01100001101111100111011,
01100001111010111000010,
01100010000101000111101,
01100010010000011000100,
01100010011011101001011,
01100010100110111010010,
01100010110010001011010,
01100010111101011100001,
01100011001000101101000,
01100011010011111101111,
01100011011111001110110,
01100011101010011111101,
01100011110101110000101,
01100011111111111111111,
01100100001011010000111,
01100100010110100001110,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000,
00000000000000000000000
);

type eg_pt_lut_array is array (0 to 2**(D_S_I_EG_V2.et_high-D_S_I_EG_V2.et_low+1)-1) of sfixed(9 downto -17);

constant EG_PT_LUT_SFIXED : eg_pt_lut_array := (
00000000001001100110011001,
00000000011001100110011001,
00000000101001100110011001,
00000000111001100110011001,
00000001001001100110011001,
00000001011001100110011001,
00000001101001100110011001,
00000001111001100110011001,
00000010001001100110011001,
00000010011001100110011001,
00000010101001100110011001,
00000010111001100110011001,
00000011001001100110011001,
00000011011001100110011001,
00000011101001100110011001,
00000011111001100110011001,
00000100001001100110011001,
00000100011001100110011001,
00000100101001100110011001,
00000100111001100110011001,
00000101001001100110011001,
00000101011001100110011001,
00000101101001100110011001,
00000101111001100110011001,
00000110001001100110011001,
00000110011001100110011001,
00000110101001100110011001,
00000110111001100110011001,
00000111001001100110011001,
00000111011001100110011001,
00000111101001100110011001,
00000111111001100110011001,
00001000001001100110011001,
00001000011001100110011001,
00001000101001100110011001,
00001000111001100110011001,
00001001001001100110011001,
00001001011001100110011001,
00001001101001100110011001,
00001001111001100110011001,
00001010001001100110011001,
00001010011001100110011001,
00001010101001100110011001,
00001010111001100110011001,
00001011001001100110011001,
00001011011001100110011001,
00001011101001100110011001,
00001011111001100110011001,
00001100001001100110011001,
00001100011001100110011001,
00001100101001100110011001,
00001100111001100110011001,
00001101001001100110011001,
00001101011001100110011001,
00001101101001100110011001,
00001101111001100110011001,
00001110001001100110011001,
00001110011001100110011001,
00001110101001100110011001,
00001110111001100110011001,
00001111001001100110011001,
00001111011001100110011001,
00001111101001100110011001,
00001111111001100110011001,
00010000001001100110011001,
00010000011001100110011001,
00010000101001100110011001,
00010000111001100110011001,
00010001001001100110011001,
00010001011001100110011001,
00010001101001100110011001,
00010001111001100110011001,
00010010001001100110011001,
00010010011001100110011001,
00010010101001100110011001,
00010010111001100110011001,
00010011001001100110011001,
00010011011001100110011001,
00010011101001100110011001,
00010011111001100110011001,
00010100001001100110011001,
00010100011001100110011001,
00010100101001100110011001,
00010100111001100110011001,
00010101001001100110011001,
00010101011001100110011001,
00010101101001100110011001,
00010101111001100110011001,
00010110001001100110011001,
00010110011001100110011001,
00010110101001100110011001,
00010110111001100110011001,
00010111001001100110011001,
00010111011001100110011001,
00010111101001100110011001,
00010111111001100110011001,
00011000001001100110011001,
00011000011001100110011001,
00011000101001100110011001,
00011000111001100110011001,
00011001001001100110011001,
00011001011001100110011001,
00011001101001100110011001,
00011001111001100110011001,
00011010001001100110011001,
00011010011001100110011001,
00011010101001100110011001,
00011010111001100110011001,
00011011001001100110011001,
00011011011001100110011001,
00011011101001100110011001,
00011011111001100110011001,
00011100001001100110011001,
00011100011001100110011001,
00011100101001100110011001,
00011100111001100110011001,
00011101001001100110011001,
00011101011001100110011001,
00011101101001100110011001,
00011101111001100110011001,
00011110001001100110011001,
00011110011001100110011001,
00011110101001100110011001,
00011110111001100110011001,
00011111001001100110011001,
00011111011001100110011001,
00011111101001100110011001,
00011111111001100110011001,
00100000001001100110011001,
00100000011001100110011001,
00100000101001100110011001,
00100000111001100110011001,
00100001001001100110011001,
00100001011001100110011001,
00100001101001100110011001,
00100001111001100110011001,
00100010001001100110011001,
00100010011001100110011001,
00100010101001100110011001,
00100010111001100110011001,
00100011001001100110011001,
00100011011001100110011001,
00100011101001100110011001,
00100011111001100110011001,
00100100001001100110011001,
00100100011001100110011001,
00100100101001100110011001,
00100100111001100110011001,
00100101001001100110011001,
00100101011001100110011001,
00100101101001100110011001,
00100101111001100110011001,
00100110001001100110011001,
00100110011001100110011001,
00100110101001100110011001,
00100110111001100110011001,
00100111001001100110011001,
00100111011001100110011001,
00100111101001100110011001,
00100111111001100110011001,
00101000001001100110011001,
00101000011001100110011001,
00101000101001100110011001,
00101000111001100110011001,
00101001001001100110011001,
00101001011001100110011001,
00101001101001100110011001,
00101001111001100110011001,
00101010001001100110011001,
00101010011001100110011001,
00101010101001100110011001,
00101010111001100110011001,
00101011001001100110011001,
00101011011001100110011001,
00101011101001100110011001,
00101011111001100110011001,
00101100001001100110011001,
00101100011001100110011001,
00101100101001100110011001,
00101100111001100110011001,
00101101001001100110011001,
00101101011001100110011001,
00101101101001100110011001,
00101101111001100110011001,
00101110001001100110011001,
00101110011001100110011001,
00101110101001100110011001,
00101110111001100110011001,
00101111001001100110011001,
00101111011001100110011001,
00101111101001100110011001,
00101111111001100110011001,
00110000001001100110011001,
00110000011001100110011001,
00110000101001100110011001,
00110000111001100110011001,
00110001001001100110011001,
00110001011001100110011001,
00110001101001100110011001,
00110001111001100110011001,
00110010001001100110011001,
00110010011001100110011001,
00110010101001100110011001,
00110010111001100110011001,
00110011001001100110011001,
00110011011001100110011001,
00110011101001100110011001,
00110011111001100110011001,
00110100001001100110011001,
00110100011001100110011001,
00110100101001100110011001,
00110100111001100110011001,
00110101001001100110011001,
00110101011001100110011001,
00110101101001100110011001,
00110101111001100110011001,
00110110001001100110011001,
00110110011001100110011001,
00110110101001100110011001,
00110110111001100110011001,
00110111001001100110011001,
00110111011001100110011001,
00110111101001100110011001,
00110111111001100110011001,
00111000001001100110011001,
00111000011001100110011001,
00111000101001100110011001,
00111000111001100110011001,
00111001001001100110011001,
00111001011001100110011001,
00111001101001100110011001,
00111001111001100110011001,
00111010001001100110011001,
00111010011001100110011001,
00111010101001100110011001,
00111010111001100110011001,
00111011001001100110011001,
00111011011001100110011001,
00111011101001100110011001,
00111011111001100110011001,
00111100001001100110011001,
00111100011001100110011001,
00111100101001100110011001,
00111100111001100110011001,
00111101001001100110011001,
00111101011001100110011001,
00111101101001100110011001,
00111101111001100110011001,
00111110001001100110011001,
00111110011001100110011001,
00111110101001100110011001,
00111110111001100110011001,
00111111001001100110011001,
00111111011001100110011001,
00111111101001100110011001,
00111111111001100110011001,
01000000001001100110011001,
01000000011001100110011001,
01000000101001100110011001,
01000000111001100110011001,
01000001001001100110011001,
01000001011001100110011001,
01000001101001100110011001,
01000001111001100110011001,
01000010001001100110011001,
01000010011001100110011001,
01000010101001100110011001,
01000010111001100110011001,
01000011001001100110011001,
01000011011001100110011001,
01000011101001100110011001,
01000011111001100110011001,
01000100001001100110011001,
01000100011001100110011001,
01000100101001100110011001,
01000100111001100110011001,
01000101001001100110011001,
01000101011001100110011001,
01000101101001100110011001,
01000101111001100110011001,
01000110001001100110011001,
01000110011001100110011001,
01000110101001100110011001,
01000110111001100110011001,
01000111001001100110011001,
01000111011001100110011001,
01000111101001100110011001,
01000111111001100110011001,
01001000001001100110011001,
01001000011001100110011001,
01001000101001100110011001,
01001000111001100110011001,
01001001001001100110011001,
01001001011001100110011001,
01001001101001100110011001,
01001001111001100110011001,
01001010001001100110011001,
01001010011001100110011001,
01001010101001100110011001,
01001010111001100110011001,
01001011001001100110011001,
01001011011001100110011001,
01001011101001100110011001,
01001011111001100110011001,
01001100001001100110011001,
01001100011001100110011001,
01001100101001100110011001,
01001100111001100110011001,
01001101001001100110011001,
01001101011001100110011001,
01001101101001100110011001,
01001101111001100110011001,
01001110001001100110011001,
01001110011001100110011001,
01001110101001100110011001,
01001110111001100110011001,
01001111001001100110011001,
01001111011001100110011001,
01001111101001100110011001,
01001111111001100110011001,
01010000001001100110011001,
01010000011001100110011001,
01010000101001100110011001,
01010000111001100110011001,
01010001001001100110011001,
01010001011001100110011001,
01010001101001100110011001,
01010001111001100110011001,
01010010001001100110011001,
01010010011001100110011001,
01010010101001100110011001,
01010010111001100110011001,
01010011001001100110011001,
01010011011001100110011001,
01010011101001100110011001,
01010011111001100110011001,
01010100001001100110011001,
01010100011001100110011001,
01010100101001100110011001,
01010100111001100110011001,
01010101001001100110011001,
01010101011001100110011001,
01010101101001100110011001,
01010101111001100110011001,
01010110001001100110011001,
01010110011001100110011001,
01010110101001100110011001,
01010110111001100110011001,
01010111001001100110011001,
01010111011001100110011001,
01010111101001100110011001,
01010111111001100110011001,
01011000001001100110011001,
01011000011001100110011001,
01011000101001100110011001,
01011000111001100110011001,
01011001001001100110011001,
01011001011001100110011001,
01011001101001100110011001,
01011001111001100110011001,
01011010001001100110011001,
01011010011001100110011001,
01011010101001100110011001,
01011010111001100110011001,
01011011001001100110011001,
01011011011001100110011001,
01011011101001100110011001,
01011011111001100110011001,
01011100001001100110011001,
01011100011001100110011001,
01011100101001100110011001,
01011100111001100110011001,
01011101001001100110011001,
01011101011001100110011001,
01011101101001100110011001,
01011101111001100110011001,
01011110001001100110011001,
01011110011001100110011001,
01011110101001100110011001,
01011110111001100110011001,
01011111001001100110011001,
01011111011001100110011001,
01011111101001100110011001,
01011111111001100110011001,
01100000001001100110011001,
01100000011001100110011001,
01100000101001100110011001,
01100000111001100110011001,
01100001001001100110011001,
01100001011001100110011001,
01100001101001100110011001,
01100001111001100110011001,
01100010001001100110011001,
01100010011001100110011001,
01100010101001100110011001,
01100010111001100110011001,
01100011001001100110011001,
01100011011001100110011001,
01100011101001100110011001,
01100011111001100110011001,
01100100001001100110011001,
01100100011001100110011001,
01100100101001100110011001,
01100100111001100110011001,
01100101001001100110011001,
01100101011001100110011001,
01100101101001100110011001,
01100101111001100110011001,
01100110001001100110011001,
01100110011001100110011001,
01100110101001100110011001,
01100110111001100110011001,
01100111001001100110011001,
01100111011001100110011001,
01100111101001100110011001,
01100111111001100110011001,
01101000001001100110011001,
01101000011001100110011001,
01101000101001100110011001,
01101000111001100110011001,
01101001001001100110011001,
01101001011001100110011001,
01101001101001100110011001,
01101001111001100110011001,
01101010001001100110011001,
01101010011001100110011001,
01101010101001100110011001,
01101010111001100110011001,
01101011001001100110011001,
01101011011001100110011001,
01101011101001100110011001,
01101011111001100110011001,
01101100001001100110011001,
01101100011001100110011001,
01101100101001100110011001,
01101100111001100110011001,
01101101001001100110011001,
01101101011001100110011001,
01101101101001100110011001,
01101101111001100110011001,
01101110001001100110011001,
01101110011001100110011001,
01101110101001100110011001,
01101110111001100110011001,
01101111001001100110011001,
01101111011001100110011001,
01101111101001100110011001,
01101111111001100110011001,
01110000001001100110011001,
01110000011001100110011001,
01110000101001100110011001,
01110000111001100110011001,
01110001001001100110011001,
01110001011001100110011001,
01110001101001100110011001,
01110001111001100110011001,
01110010001001100110011001,
01110010011001100110011001,
01110010101001100110011001,
01110010111001100110011001,
01110011001001100110011001,
01110011011001100110011001,
01110011101001100110011001,
01110011111001100110011001,
01110100001001100110011001,
01110100011001100110011001,
01110100101001100110011001,
01110100111001100110011001,
01110101001001100110011001,
01110101011001100110011001,
01110101101001100110011001,
01110101111001100110011001,
01110110001001100110011001,
01110110011001100110011001,
01110110101001100110011001,
01110110111001100110011001,
01110111001001100110011001,
01110111011001100110011001,
01110111101001100110011001,
01110111111001100110011001,
01111000001001100110011001,
01111000011001100110011001,
01111000101001100110011001,
01111000111001100110011001,
01111001001001100110011001,
01111001011001100110011001,
01111001101001100110011001,
01111001111001100110011001,
01111010001001100110011001,
01111010011001100110011001,
01111010101001100110011001,
01111010111001100110011001,
01111011001001100110011001,
01111011011001100110011001,
01111011101001100110011001,
01111011111001100110011001,
01111100001001100110011001,
01111100011001100110011001,
01111100101001100110011001,
01111100111001100110011001,
01111101001001100110011001,
01111101011001100110011001,
01111101101001100110011001,
01111101111001100110011001,
01111110001001100110011001,
01111110011001100110011001,
01111110101001100110011001,
01111110111001100110011001,
01111111001001100110011001,
01111111011001100110011001,
01111111101001100110011001,
01111111111001100110011001
);

constant TAU_PT_LUT_SFIXED : eg_pt_lut_array := EG_PT_LUT_SFIXED;

type jet_pt_lut_array is array (0 to 2**(D_S_I_JET_V2.et_high-D_S_I_JET_V2.et_low+1)-1) of sfixed(11 downto -17);

constant JET_PT_LUT_SFIXED : jet_pt_lut_array := (
0000000000001001100110011001,
0000000000011001100110011001,
0000000000101001100110011001,
0000000000111001100110011001,
0000000001001001100110011001,
0000000001011001100110011001,
0000000001101001100110011001,
0000000001111001100110011001,
0000000010001001100110011001,
0000000010011001100110011001,
0000000010101001100110011001,
0000000010111001100110011001,
0000000011001001100110011001,
0000000011011001100110011001,
0000000011101001100110011001,
0000000011111001100110011001,
0000000100001001100110011001,
0000000100011001100110011001,
0000000100101001100110011001,
0000000100111001100110011001,
0000000101001001100110011001,
0000000101011001100110011001,
0000000101101001100110011001,
0000000101111001100110011001,
0000000110001001100110011001,
0000000110011001100110011001,
0000000110101001100110011001,
0000000110111001100110011001,
0000000111001001100110011001,
0000000111011001100110011001,
0000000111101001100110011001,
0000000111111001100110011001,
0000001000001001100110011001,
0000001000011001100110011001,
0000001000101001100110011001,
0000001000111001100110011001,
0000001001001001100110011001,
0000001001011001100110011001,
0000001001101001100110011001,
0000001001111001100110011001,
0000001010001001100110011001,
0000001010011001100110011001,
0000001010101001100110011001,
0000001010111001100110011001,
0000001011001001100110011001,
0000001011011001100110011001,
0000001011101001100110011001,
0000001011111001100110011001,
0000001100001001100110011001,
0000001100011001100110011001,
0000001100101001100110011001,
0000001100111001100110011001,
0000001101001001100110011001,
0000001101011001100110011001,
0000001101101001100110011001,
0000001101111001100110011001,
0000001110001001100110011001,
0000001110011001100110011001,
0000001110101001100110011001,
0000001110111001100110011001,
0000001111001001100110011001,
0000001111011001100110011001,
0000001111101001100110011001,
0000001111111001100110011001,
0000010000001001100110011001,
0000010000011001100110011001,
0000010000101001100110011001,
0000010000111001100110011001,
0000010001001001100110011001,
0000010001011001100110011001,
0000010001101001100110011001,
0000010001111001100110011001,
0000010010001001100110011001,
0000010010011001100110011001,
0000010010101001100110011001,
0000010010111001100110011001,
0000010011001001100110011001,
0000010011011001100110011001,
0000010011101001100110011001,
0000010011111001100110011001,
0000010100001001100110011001,
0000010100011001100110011001,
0000010100101001100110011001,
0000010100111001100110011001,
0000010101001001100110011001,
0000010101011001100110011001,
0000010101101001100110011001,
0000010101111001100110011001,
0000010110001001100110011001,
0000010110011001100110011001,
0000010110101001100110011001,
0000010110111001100110011001,
0000010111001001100110011001,
0000010111011001100110011001,
0000010111101001100110011001,
0000010111111001100110011001,
0000011000001001100110011001,
0000011000011001100110011001,
0000011000101001100110011001,
0000011000111001100110011001,
0000011001001001100110011001,
0000011001011001100110011001,
0000011001101001100110011001,
0000011001111001100110011001,
0000011010001001100110011001,
0000011010011001100110011001,
0000011010101001100110011001,
0000011010111001100110011001,
0000011011001001100110011001,
0000011011011001100110011001,
0000011011101001100110011001,
0000011011111001100110011001,
0000011100001001100110011001,
0000011100011001100110011001,
0000011100101001100110011001,
0000011100111001100110011001,
0000011101001001100110011001,
0000011101011001100110011001,
0000011101101001100110011001,
0000011101111001100110011001,
0000011110001001100110011001,
0000011110011001100110011001,
0000011110101001100110011001,
0000011110111001100110011001,
0000011111001001100110011001,
0000011111011001100110011001,
0000011111101001100110011001,
0000011111111001100110011001,
0000100000001001100110011001,
0000100000011001100110011001,
0000100000101001100110011001,
0000100000111001100110011001,
0000100001001001100110011001,
0000100001011001100110011001,
0000100001101001100110011001,
0000100001111001100110011001,
0000100010001001100110011001,
0000100010011001100110011001,
0000100010101001100110011001,
0000100010111001100110011001,
0000100011001001100110011001,
0000100011011001100110011001,
0000100011101001100110011001,
0000100011111001100110011001,
0000100100001001100110011001,
0000100100011001100110011001,
0000100100101001100110011001,
0000100100111001100110011001,
0000100101001001100110011001,
0000100101011001100110011001,
0000100101101001100110011001,
0000100101111001100110011001,
0000100110001001100110011001,
0000100110011001100110011001,
0000100110101001100110011001,
0000100110111001100110011001,
0000100111001001100110011001,
0000100111011001100110011001,
0000100111101001100110011001,
0000100111111001100110011001,
0000101000001001100110011001,
0000101000011001100110011001,
0000101000101001100110011001,
0000101000111001100110011001,
0000101001001001100110011001,
0000101001011001100110011001,
0000101001101001100110011001,
0000101001111001100110011001,
0000101010001001100110011001,
0000101010011001100110011001,
0000101010101001100110011001,
0000101010111001100110011001,
0000101011001001100110011001,
0000101011011001100110011001,
0000101011101001100110011001,
0000101011111001100110011001,
0000101100001001100110011001,
0000101100011001100110011001,
0000101100101001100110011001,
0000101100111001100110011001,
0000101101001001100110011001,
0000101101011001100110011001,
0000101101101001100110011001,
0000101101111001100110011001,
0000101110001001100110011001,
0000101110011001100110011001,
0000101110101001100110011001,
0000101110111001100110011001,
0000101111001001100110011001,
0000101111011001100110011001,
0000101111101001100110011001,
0000101111111001100110011001,
0000110000001001100110011001,
0000110000011001100110011001,
0000110000101001100110011001,
0000110000111001100110011001,
0000110001001001100110011001,
0000110001011001100110011001,
0000110001101001100110011001,
0000110001111001100110011001,
0000110010001001100110011001,
0000110010011001100110011001,
0000110010101001100110011001,
0000110010111001100110011001,
0000110011001001100110011001,
0000110011011001100110011001,
0000110011101001100110011001,
0000110011111001100110011001,
0000110100001001100110011001,
0000110100011001100110011001,
0000110100101001100110011001,
0000110100111001100110011001,
0000110101001001100110011001,
0000110101011001100110011001,
0000110101101001100110011001,
0000110101111001100110011001,
0000110110001001100110011001,
0000110110011001100110011001,
0000110110101001100110011001,
0000110110111001100110011001,
0000110111001001100110011001,
0000110111011001100110011001,
0000110111101001100110011001,
0000110111111001100110011001,
0000111000001001100110011001,
0000111000011001100110011001,
0000111000101001100110011001,
0000111000111001100110011001,
0000111001001001100110011001,
0000111001011001100110011001,
0000111001101001100110011001,
0000111001111001100110011001,
0000111010001001100110011001,
0000111010011001100110011001,
0000111010101001100110011001,
0000111010111001100110011001,
0000111011001001100110011001,
0000111011011001100110011001,
0000111011101001100110011001,
0000111011111001100110011001,
0000111100001001100110011001,
0000111100011001100110011001,
0000111100101001100110011001,
0000111100111001100110011001,
0000111101001001100110011001,
0000111101011001100110011001,
0000111101101001100110011001,
0000111101111001100110011001,
0000111110001001100110011001,
0000111110011001100110011001,
0000111110101001100110011001,
0000111110111001100110011001,
0000111111001001100110011001,
0000111111011001100110011001,
0000111111101001100110011001,
0000111111111001100110011001,
0001000000001001100110011001,
0001000000011001100110011001,
0001000000101001100110011001,
0001000000111001100110011001,
0001000001001001100110011001,
0001000001011001100110011001,
0001000001101001100110011001,
0001000001111001100110011001,
0001000010001001100110011001,
0001000010011001100110011001,
0001000010101001100110011001,
0001000010111001100110011001,
0001000011001001100110011001,
0001000011011001100110011001,
0001000011101001100110011001,
0001000011111001100110011001,
0001000100001001100110011001,
0001000100011001100110011001,
0001000100101001100110011001,
0001000100111001100110011001,
0001000101001001100110011001,
0001000101011001100110011001,
0001000101101001100110011001,
0001000101111001100110011001,
0001000110001001100110011001,
0001000110011001100110011001,
0001000110101001100110011001,
0001000110111001100110011001,
0001000111001001100110011001,
0001000111011001100110011001,
0001000111101001100110011001,
0001000111111001100110011001,
0001001000001001100110011001,
0001001000011001100110011001,
0001001000101001100110011001,
0001001000111001100110011001,
0001001001001001100110011001,
0001001001011001100110011001,
0001001001101001100110011001,
0001001001111001100110011001,
0001001010001001100110011001,
0001001010011001100110011001,
0001001010101001100110011001,
0001001010111001100110011001,
0001001011001001100110011001,
0001001011011001100110011001,
0001001011101001100110011001,
0001001011111001100110011001,
0001001100001001100110011001,
0001001100011001100110011001,
0001001100101001100110011001,
0001001100111001100110011001,
0001001101001001100110011001,
0001001101011001100110011001,
0001001101101001100110011001,
0001001101111001100110011001,
0001001110001001100110011001,
0001001110011001100110011001,
0001001110101001100110011001,
0001001110111001100110011001,
0001001111001001100110011001,
0001001111011001100110011001,
0001001111101001100110011001,
0001001111111001100110011001,
0001010000001001100110011001,
0001010000011001100110011001,
0001010000101001100110011001,
0001010000111001100110011001,
0001010001001001100110011001,
0001010001011001100110011001,
0001010001101001100110011001,
0001010001111001100110011001,
0001010010001001100110011001,
0001010010011001100110011001,
0001010010101001100110011001,
0001010010111001100110011001,
0001010011001001100110011001,
0001010011011001100110011001,
0001010011101001100110011001,
0001010011111001100110011001,
0001010100001001100110011001,
0001010100011001100110011001,
0001010100101001100110011001,
0001010100111001100110011001,
0001010101001001100110011001,
0001010101011001100110011001,
0001010101101001100110011001,
0001010101111001100110011001,
0001010110001001100110011001,
0001010110011001100110011001,
0001010110101001100110011001,
0001010110111001100110011001,
0001010111001001100110011001,
0001010111011001100110011001,
0001010111101001100110011001,
0001010111111001100110011001,
0001011000001001100110011001,
0001011000011001100110011001,
0001011000101001100110011001,
0001011000111001100110011001,
0001011001001001100110011001,
0001011001011001100110011001,
0001011001101001100110011001,
0001011001111001100110011001,
0001011010001001100110011001,
0001011010011001100110011001,
0001011010101001100110011001,
0001011010111001100110011001,
0001011011001001100110011001,
0001011011011001100110011001,
0001011011101001100110011001,
0001011011111001100110011001,
0001011100001001100110011001,
0001011100011001100110011001,
0001011100101001100110011001,
0001011100111001100110011001,
0001011101001001100110011001,
0001011101011001100110011001,
0001011101101001100110011001,
0001011101111001100110011001,
0001011110001001100110011001,
0001011110011001100110011001,
0001011110101001100110011001,
0001011110111001100110011001,
0001011111001001100110011001,
0001011111011001100110011001,
0001011111101001100110011001,
0001011111111001100110011001,
0001100000001001100110011001,
0001100000011001100110011001,
0001100000101001100110011001,
0001100000111001100110011001,
0001100001001001100110011001,
0001100001011001100110011001,
0001100001101001100110011001,
0001100001111001100110011001,
0001100010001001100110011001,
0001100010011001100110011001,
0001100010101001100110011001,
0001100010111001100110011001,
0001100011001001100110011001,
0001100011011001100110011001,
0001100011101001100110011001,
0001100011111001100110011001,
0001100100001001100110011001,
0001100100011001100110011001,
0001100100101001100110011001,
0001100100111001100110011001,
0001100101001001100110011001,
0001100101011001100110011001,
0001100101101001100110011001,
0001100101111001100110011001,
0001100110001001100110011001,
0001100110011001100110011001,
0001100110101001100110011001,
0001100110111001100110011001,
0001100111001001100110011001,
0001100111011001100110011001,
0001100111101001100110011001,
0001100111111001100110011001,
0001101000001001100110011001,
0001101000011001100110011001,
0001101000101001100110011001,
0001101000111001100110011001,
0001101001001001100110011001,
0001101001011001100110011001,
0001101001101001100110011001,
0001101001111001100110011001,
0001101010001001100110011001,
0001101010011001100110011001,
0001101010101001100110011001,
0001101010111001100110011001,
0001101011001001100110011001,
0001101011011001100110011001,
0001101011101001100110011001,
0001101011111001100110011001,
0001101100001001100110011001,
0001101100011001100110011001,
0001101100101001100110011001,
0001101100111001100110011001,
0001101101001001100110011001,
0001101101011001100110011001,
0001101101101001100110011001,
0001101101111001100110011001,
0001101110001001100110011001,
0001101110011001100110011001,
0001101110101001100110011001,
0001101110111001100110011001,
0001101111001001100110011001,
0001101111011001100110011001,
0001101111101001100110011001,
0001101111111001100110011001,
0001110000001001100110011001,
0001110000011001100110011001,
0001110000101001100110011001,
0001110000111001100110011001,
0001110001001001100110011001,
0001110001011001100110011001,
0001110001101001100110011001,
0001110001111001100110011001,
0001110010001001100110011001,
0001110010011001100110011001,
0001110010101001100110011001,
0001110010111001100110011001,
0001110011001001100110011001,
0001110011011001100110011001,
0001110011101001100110011001,
0001110011111001100110011001,
0001110100001001100110011001,
0001110100011001100110011001,
0001110100101001100110011001,
0001110100111001100110011001,
0001110101001001100110011001,
0001110101011001100110011001,
0001110101101001100110011001,
0001110101111001100110011001,
0001110110001001100110011001,
0001110110011001100110011001,
0001110110101001100110011001,
0001110110111001100110011001,
0001110111001001100110011001,
0001110111011001100110011001,
0001110111101001100110011001,
0001110111111001100110011001,
0001111000001001100110011001,
0001111000011001100110011001,
0001111000101001100110011001,
0001111000111001100110011001,
0001111001001001100110011001,
0001111001011001100110011001,
0001111001101001100110011001,
0001111001111001100110011001,
0001111010001001100110011001,
0001111010011001100110011001,
0001111010101001100110011001,
0001111010111001100110011001,
0001111011001001100110011001,
0001111011011001100110011001,
0001111011101001100110011001,
0001111011111001100110011001,
0001111100001001100110011001,
0001111100011001100110011001,
0001111100101001100110011001,
0001111100111001100110011001,
0001111101001001100110011001,
0001111101011001100110011001,
0001111101101001100110011001,
0001111101111001100110011001,
0001111110001001100110011001,
0001111110011001100110011001,
0001111110101001100110011001,
0001111110111001100110011001,
0001111111001001100110011001,
0001111111011001100110011001,
0001111111101001100110011001,
0001111111111001100110011001,
0010000000001001100110011001,
0010000000011001100110011001,
0010000000101001100110011001,
0010000000111001100110011001,
0010000001001001100110011001,
0010000001011001100110011001,
0010000001101001100110011001,
0010000001111001100110011001,
0010000010001001100110011001,
0010000010011001100110011001,
0010000010101001100110011001,
0010000010111001100110011001,
0010000011001001100110011001,
0010000011011001100110011001,
0010000011101001100110011001,
0010000011111001100110011001,
0010000100001001100110011001,
0010000100011001100110011001,
0010000100101001100110011001,
0010000100111001100110011001,
0010000101001001100110011001,
0010000101011001100110011001,
0010000101101001100110011001,
0010000101111001100110011001,
0010000110001001100110011001,
0010000110011001100110011001,
0010000110101001100110011001,
0010000110111001100110011001,
0010000111001001100110011001,
0010000111011001100110011001,
0010000111101001100110011001,
0010000111111001100110011001,
0010001000001001100110011001,
0010001000011001100110011001,
0010001000101001100110011001,
0010001000111001100110011001,
0010001001001001100110011001,
0010001001011001100110011001,
0010001001101001100110011001,
0010001001111001100110011001,
0010001010001001100110011001,
0010001010011001100110011001,
0010001010101001100110011001,
0010001010111001100110011001,
0010001011001001100110011001,
0010001011011001100110011001,
0010001011101001100110011001,
0010001011111001100110011001,
0010001100001001100110011001,
0010001100011001100110011001,
0010001100101001100110011001,
0010001100111001100110011001,
0010001101001001100110011001,
0010001101011001100110011001,
0010001101101001100110011001,
0010001101111001100110011001,
0010001110001001100110011001,
0010001110011001100110011001,
0010001110101001100110011001,
0010001110111001100110011001,
0010001111001001100110011001,
0010001111011001100110011001,
0010001111101001100110011001,
0010001111111001100110011001,
0010010000001001100110011001,
0010010000011001100110011001,
0010010000101001100110011001,
0010010000111001100110011001,
0010010001001001100110011001,
0010010001011001100110011001,
0010010001101001100110011001,
0010010001111001100110011001,
0010010010001001100110011001,
0010010010011001100110011001,
0010010010101001100110011001,
0010010010111001100110011001,
0010010011001001100110011001,
0010010011011001100110011001,
0010010011101001100110011001,
0010010011111001100110011001,
0010010100001001100110011001,
0010010100011001100110011001,
0010010100101001100110011001,
0010010100111001100110011001,
0010010101001001100110011001,
0010010101011001100110011001,
0010010101101001100110011001,
0010010101111001100110011001,
0010010110001001100110011001,
0010010110011001100110011001,
0010010110101001100110011001,
0010010110111001100110011001,
0010010111001001100110011001,
0010010111011001100110011001,
0010010111101001100110011001,
0010010111111001100110011001,
0010011000001001100110011001,
0010011000011001100110011001,
0010011000101001100110011001,
0010011000111001100110011001,
0010011001001001100110011001,
0010011001011001100110011001,
0010011001101001100110011001,
0010011001111001100110011001,
0010011010001001100110011001,
0010011010011001100110011001,
0010011010101001100110011001,
0010011010111001100110011001,
0010011011001001100110011001,
0010011011011001100110011001,
0010011011101001100110011001,
0010011011111001100110011001,
0010011100001001100110011001,
0010011100011001100110011001,
0010011100101001100110011001,
0010011100111001100110011001,
0010011101001001100110011001,
0010011101011001100110011001,
0010011101101001100110011001,
0010011101111001100110011001,
0010011110001001100110011001,
0010011110011001100110011001,
0010011110101001100110011001,
0010011110111001100110011001,
0010011111001001100110011001,
0010011111011001100110011001,
0010011111101001100110011001,
0010011111111001100110011001,
0010100000001001100110011001,
0010100000011001100110011001,
0010100000101001100110011001,
0010100000111001100110011001,
0010100001001001100110011001,
0010100001011001100110011001,
0010100001101001100110011001,
0010100001111001100110011001,
0010100010001001100110011001,
0010100010011001100110011001,
0010100010101001100110011001,
0010100010111001100110011001,
0010100011001001100110011001,
0010100011011001100110011001,
0010100011101001100110011001,
0010100011111001100110011001,
0010100100001001100110011001,
0010100100011001100110011001,
0010100100101001100110011001,
0010100100111001100110011001,
0010100101001001100110011001,
0010100101011001100110011001,
0010100101101001100110011001,
0010100101111001100110011001,
0010100110001001100110011001,
0010100110011001100110011001,
0010100110101001100110011001,
0010100110111001100110011001,
0010100111001001100110011001,
0010100111011001100110011001,
0010100111101001100110011001,
0010100111111001100110011001,
0010101000001001100110011001,
0010101000011001100110011001,
0010101000101001100110011001,
0010101000111001100110011001,
0010101001001001100110011001,
0010101001011001100110011001,
0010101001101001100110011001,
0010101001111001100110011001,
0010101010001001100110011001,
0010101010011001100110011001,
0010101010101001100110011001,
0010101010111001100110011001,
0010101011001001100110011001,
0010101011011001100110011001,
0010101011101001100110011001,
0010101011111001100110011001,
0010101100001001100110011001,
0010101100011001100110011001,
0010101100101001100110011001,
0010101100111001100110011001,
0010101101001001100110011001,
0010101101011001100110011001,
0010101101101001100110011001,
0010101101111001100110011001,
0010101110001001100110011001,
0010101110011001100110011001,
0010101110101001100110011001,
0010101110111001100110011001,
0010101111001001100110011001,
0010101111011001100110011001,
0010101111101001100110011001,
0010101111111001100110011001,
0010110000001001100110011001,
0010110000011001100110011001,
0010110000101001100110011001,
0010110000111001100110011001,
0010110001001001100110011001,
0010110001011001100110011001,
0010110001101001100110011001,
0010110001111001100110011001,
0010110010001001100110011001,
0010110010011001100110011001,
0010110010101001100110011001,
0010110010111001100110011001,
0010110011001001100110011001,
0010110011011001100110011001,
0010110011101001100110011001,
0010110011111001100110011001,
0010110100001001100110011001,
0010110100011001100110011001,
0010110100101001100110011001,
0010110100111001100110011001,
0010110101001001100110011001,
0010110101011001100110011001,
0010110101101001100110011001,
0010110101111001100110011001,
0010110110001001100110011001,
0010110110011001100110011001,
0010110110101001100110011001,
0010110110111001100110011001,
0010110111001001100110011001,
0010110111011001100110011001,
0010110111101001100110011001,
0010110111111001100110011001,
0010111000001001100110011001,
0010111000011001100110011001,
0010111000101001100110011001,
0010111000111001100110011001,
0010111001001001100110011001,
0010111001011001100110011001,
0010111001101001100110011001,
0010111001111001100110011001,
0010111010001001100110011001,
0010111010011001100110011001,
0010111010101001100110011001,
0010111010111001100110011001,
0010111011001001100110011001,
0010111011011001100110011001,
0010111011101001100110011001,
0010111011111001100110011001,
0010111100001001100110011001,
0010111100011001100110011001,
0010111100101001100110011001,
0010111100111001100110011001,
0010111101001001100110011001,
0010111101011001100110011001,
0010111101101001100110011001,
0010111101111001100110011001,
0010111110001001100110011001,
0010111110011001100110011001,
0010111110101001100110011001,
0010111110111001100110011001,
0010111111001001100110011001,
0010111111011001100110011001,
0010111111101001100110011001,
0010111111111001100110011001,
0011000000001001100110011001,
0011000000011001100110011001,
0011000000101001100110011001,
0011000000111001100110011001,
0011000001001001100110011001,
0011000001011001100110011001,
0011000001101001100110011001,
0011000001111001100110011001,
0011000010001001100110011001,
0011000010011001100110011001,
0011000010101001100110011001,
0011000010111001100110011001,
0011000011001001100110011001,
0011000011011001100110011001,
0011000011101001100110011001,
0011000011111001100110011001,
0011000100001001100110011001,
0011000100011001100110011001,
0011000100101001100110011001,
0011000100111001100110011001,
0011000101001001100110011001,
0011000101011001100110011001,
0011000101101001100110011001,
0011000101111001100110011001,
0011000110001001100110011001,
0011000110011001100110011001,
0011000110101001100110011001,
0011000110111001100110011001,
0011000111001001100110011001,
0011000111011001100110011001,
0011000111101001100110011001,
0011000111111001100110011001,
0011001000001001100110011001,
0011001000011001100110011001,
0011001000101001100110011001,
0011001000111001100110011001,
0011001001001001100110011001,
0011001001011001100110011001,
0011001001101001100110011001,
0011001001111001100110011001,
0011001010001001100110011001,
0011001010011001100110011001,
0011001010101001100110011001,
0011001010111001100110011001,
0011001011001001100110011001,
0011001011011001100110011001,
0011001011101001100110011001,
0011001011111001100110011001,
0011001100001001100110011001,
0011001100011001100110011001,
0011001100101001100110011001,
0011001100111001100110011001,
0011001101001001100110011001,
0011001101011001100110011001,
0011001101101001100110011001,
0011001101111001100110011001,
0011001110001001100110011001,
0011001110011001100110011001,
0011001110101001100110011001,
0011001110111001100110011001,
0011001111001001100110011001,
0011001111011001100110011001,
0011001111101001100110011001,
0011001111111001100110011001,
0011010000001001100110011001,
0011010000011001100110011001,
0011010000101001100110011001,
0011010000111001100110011001,
0011010001001001100110011001,
0011010001011001100110011001,
0011010001101001100110011001,
0011010001111001100110011001,
0011010010001001100110011001,
0011010010011001100110011001,
0011010010101001100110011001,
0011010010111001100110011001,
0011010011001001100110011001,
0011010011011001100110011001,
0011010011101001100110011001,
0011010011111001100110011001,
0011010100001001100110011001,
0011010100011001100110011001,
0011010100101001100110011001,
0011010100111001100110011001,
0011010101001001100110011001,
0011010101011001100110011001,
0011010101101001100110011001,
0011010101111001100110011001,
0011010110001001100110011001,
0011010110011001100110011001,
0011010110101001100110011001,
0011010110111001100110011001,
0011010111001001100110011001,
0011010111011001100110011001,
0011010111101001100110011001,
0011010111111001100110011001,
0011011000001001100110011001,
0011011000011001100110011001,
0011011000101001100110011001,
0011011000111001100110011001,
0011011001001001100110011001,
0011011001011001100110011001,
0011011001101001100110011001,
0011011001111001100110011001,
0011011010001001100110011001,
0011011010011001100110011001,
0011011010101001100110011001,
0011011010111001100110011001,
0011011011001001100110011001,
0011011011011001100110011001,
0011011011101001100110011001,
0011011011111001100110011001,
0011011100001001100110011001,
0011011100011001100110011001,
0011011100101001100110011001,
0011011100111001100110011001,
0011011101001001100110011001,
0011011101011001100110011001,
0011011101101001100110011001,
0011011101111001100110011001,
0011011110001001100110011001,
0011011110011001100110011001,
0011011110101001100110011001,
0011011110111001100110011001,
0011011111001001100110011001,
0011011111011001100110011001,
0011011111101001100110011001,
0011011111111001100110011001,
0011100000001001100110011001,
0011100000011001100110011001,
0011100000101001100110011001,
0011100000111001100110011001,
0011100001001001100110011001,
0011100001011001100110011001,
0011100001101001100110011001,
0011100001111001100110011001,
0011100010001001100110011001,
0011100010011001100110011001,
0011100010101001100110011001,
0011100010111001100110011001,
0011100011001001100110011001,
0011100011011001100110011001,
0011100011101001100110011001,
0011100011111001100110011001,
0011100100001001100110011001,
0011100100011001100110011001,
0011100100101001100110011001,
0011100100111001100110011001,
0011100101001001100110011001,
0011100101011001100110011001,
0011100101101001100110011001,
0011100101111001100110011001,
0011100110001001100110011001,
0011100110011001100110011001,
0011100110101001100110011001,
0011100110111001100110011001,
0011100111001001100110011001,
0011100111011001100110011001,
0011100111101001100110011001,
0011100111111001100110011001,
0011101000001001100110011001,
0011101000011001100110011001,
0011101000101001100110011001,
0011101000111001100110011001,
0011101001001001100110011001,
0011101001011001100110011001,
0011101001101001100110011001,
0011101001111001100110011001,
0011101010001001100110011001,
0011101010011001100110011001,
0011101010101001100110011001,
0011101010111001100110011001,
0011101011001001100110011001,
0011101011011001100110011001,
0011101011101001100110011001,
0011101011111001100110011001,
0011101100001001100110011001,
0011101100011001100110011001,
0011101100101001100110011001,
0011101100111001100110011001,
0011101101001001100110011001,
0011101101011001100110011001,
0011101101101001100110011001,
0011101101111001100110011001,
0011101110001001100110011001,
0011101110011001100110011001,
0011101110101001100110011001,
0011101110111001100110011001,
0011101111001001100110011001,
0011101111011001100110011001,
0011101111101001100110011001,
0011101111111001100110011001,
0011110000001001100110011001,
0011110000011001100110011001,
0011110000101001100110011001,
0011110000111001100110011001,
0011110001001001100110011001,
0011110001011001100110011001,
0011110001101001100110011001,
0011110001111001100110011001,
0011110010001001100110011001,
0011110010011001100110011001,
0011110010101001100110011001,
0011110010111001100110011001,
0011110011001001100110011001,
0011110011011001100110011001,
0011110011101001100110011001,
0011110011111001100110011001,
0011110100001001100110011001,
0011110100011001100110011001,
0011110100101001100110011001,
0011110100111001100110011001,
0011110101001001100110011001,
0011110101011001100110011001,
0011110101101001100110011001,
0011110101111001100110011001,
0011110110001001100110011001,
0011110110011001100110011001,
0011110110101001100110011001,
0011110110111001100110011001,
0011110111001001100110011001,
0011110111011001100110011001,
0011110111101001100110011001,
0011110111111001100110011001,
0011111000001001100110011001,
0011111000011001100110011001,
0011111000101001100110011001,
0011111000111001100110011001,
0011111001001001100110011001,
0011111001011001100110011001,
0011111001101001100110011001,
0011111001111001100110011001,
0011111010001001100110011001,
0011111010011001100110011001,
0011111010101001100110011001,
0011111010111001100110011001,
0011111011001001100110011001,
0011111011011001100110011001,
0011111011101001100110011001,
0011111011111001100110011001,
0011111100001001100110011001,
0011111100011001100110011001,
0011111100101001100110011001,
0011111100111001100110011001,
0011111101001001100110011001,
0011111101011001100110011001,
0011111101101001100110011001,
0011111101111001100110011001,
0011111110001001100110011001,
0011111110011001100110011001,
0011111110101001100110011001,
0011111110111001100110011001,
0011111111001001100110011001,
0011111111011001100110011001,
0011111111101001100110011001,
0011111111111001100110011001,
0100000000001001100110011001,
0100000000011001100110011001,
0100000000101001100110011001,
0100000000111001100110011001,
0100000001001001100110011001,
0100000001011001100110011001,
0100000001101001100110011001,
0100000001111001100110011001,
0100000010001001100110011001,
0100000010011001100110011001,
0100000010101001100110011001,
0100000010111001100110011001,
0100000011001001100110011001,
0100000011011001100110011001,
0100000011101001100110011001,
0100000011111001100110011001,
0100000100001001100110011001,
0100000100011001100110011001,
0100000100101001100110011001,
0100000100111001100110011001,
0100000101001001100110011001,
0100000101011001100110011001,
0100000101101001100110011001,
0100000101111001100110011001,
0100000110001001100110011001,
0100000110011001100110011001,
0100000110101001100110011001,
0100000110111001100110011001,
0100000111001001100110011001,
0100000111011001100110011001,
0100000111101001100110011001,
0100000111111001100110011001,
0100001000001001100110011001,
0100001000011001100110011001,
0100001000101001100110011001,
0100001000111001100110011001,
0100001001001001100110011001,
0100001001011001100110011001,
0100001001101001100110011001,
0100001001111001100110011001,
0100001010001001100110011001,
0100001010011001100110011001,
0100001010101001100110011001,
0100001010111001100110011001,
0100001011001001100110011001,
0100001011011001100110011001,
0100001011101001100110011001,
0100001011111001100110011001,
0100001100001001100110011001,
0100001100011001100110011001,
0100001100101001100110011001,
0100001100111001100110011001,
0100001101001001100110011001,
0100001101011001100110011001,
0100001101101001100110011001,
0100001101111001100110011001,
0100001110001001100110011001,
0100001110011001100110011001,
0100001110101001100110011001,
0100001110111001100110011001,
0100001111001001100110011001,
0100001111011001100110011001,
0100001111101001100110011001,
0100001111111001100110011001,
0100010000001001100110011001,
0100010000011001100110011001,
0100010000101001100110011001,
0100010000111001100110011001,
0100010001001001100110011001,
0100010001011001100110011001,
0100010001101001100110011001,
0100010001111001100110011001,
0100010010001001100110011001,
0100010010011001100110011001,
0100010010101001100110011001,
0100010010111001100110011001,
0100010011001001100110011001,
0100010011011001100110011001,
0100010011101001100110011001,
0100010011111001100110011001,
0100010100001001100110011001,
0100010100011001100110011001,
0100010100101001100110011001,
0100010100111001100110011001,
0100010101001001100110011001,
0100010101011001100110011001,
0100010101101001100110011001,
0100010101111001100110011001,
0100010110001001100110011001,
0100010110011001100110011001,
0100010110101001100110011001,
0100010110111001100110011001,
0100010111001001100110011001,
0100010111011001100110011001,
0100010111101001100110011001,
0100010111111001100110011001,
0100011000001001100110011001,
0100011000011001100110011001,
0100011000101001100110011001,
0100011000111001100110011001,
0100011001001001100110011001,
0100011001011001100110011001,
0100011001101001100110011001,
0100011001111001100110011001,
0100011010001001100110011001,
0100011010011001100110011001,
0100011010101001100110011001,
0100011010111001100110011001,
0100011011001001100110011001,
0100011011011001100110011001,
0100011011101001100110011001,
0100011011111001100110011001,
0100011100001001100110011001,
0100011100011001100110011001,
0100011100101001100110011001,
0100011100111001100110011001,
0100011101001001100110011001,
0100011101011001100110011001,
0100011101101001100110011001,
0100011101111001100110011001,
0100011110001001100110011001,
0100011110011001100110011001,
0100011110101001100110011001,
0100011110111001100110011001,
0100011111001001100110011001,
0100011111011001100110011001,
0100011111101001100110011001,
0100011111111001100110011001,
0100100000001001100110011001,
0100100000011001100110011001,
0100100000101001100110011001,
0100100000111001100110011001,
0100100001001001100110011001,
0100100001011001100110011001,
0100100001101001100110011001,
0100100001111001100110011001,
0100100010001001100110011001,
0100100010011001100110011001,
0100100010101001100110011001,
0100100010111001100110011001,
0100100011001001100110011001,
0100100011011001100110011001,
0100100011101001100110011001,
0100100011111001100110011001,
0100100100001001100110011001,
0100100100011001100110011001,
0100100100101001100110011001,
0100100100111001100110011001,
0100100101001001100110011001,
0100100101011001100110011001,
0100100101101001100110011001,
0100100101111001100110011001,
0100100110001001100110011001,
0100100110011001100110011001,
0100100110101001100110011001,
0100100110111001100110011001,
0100100111001001100110011001,
0100100111011001100110011001,
0100100111101001100110011001,
0100100111111001100110011001,
0100101000001001100110011001,
0100101000011001100110011001,
0100101000101001100110011001,
0100101000111001100110011001,
0100101001001001100110011001,
0100101001011001100110011001,
0100101001101001100110011001,
0100101001111001100110011001,
0100101010001001100110011001,
0100101010011001100110011001,
0100101010101001100110011001,
0100101010111001100110011001,
0100101011001001100110011001,
0100101011011001100110011001,
0100101011101001100110011001,
0100101011111001100110011001,
0100101100001001100110011001,
0100101100011001100110011001,
0100101100101001100110011001,
0100101100111001100110011001,
0100101101001001100110011001,
0100101101011001100110011001,
0100101101101001100110011001,
0100101101111001100110011001,
0100101110001001100110011001,
0100101110011001100110011001,
0100101110101001100110011001,
0100101110111001100110011001,
0100101111001001100110011001,
0100101111011001100110011001,
0100101111101001100110011001,
0100101111111001100110011001,
0100110000001001100110011001,
0100110000011001100110011001,
0100110000101001100110011001,
0100110000111001100110011001,
0100110001001001100110011001,
0100110001011001100110011001,
0100110001101001100110011001,
0100110001111001100110011001,
0100110010001001100110011001,
0100110010011001100110011001,
0100110010101001100110011001,
0100110010111001100110011001,
0100110011001001100110011001,
0100110011011001100110011001,
0100110011101001100110011001,
0100110011111001100110011001,
0100110100001001100110011001,
0100110100011001100110011001,
0100110100101001100110011001,
0100110100111001100110011001,
0100110101001001100110011001,
0100110101011001100110011001,
0100110101101001100110011001,
0100110101111001100110011001,
0100110110001001100110011001,
0100110110011001100110011001,
0100110110101001100110011001,
0100110110111001100110011001,
0100110111001001100110011001,
0100110111011001100110011001,
0100110111101001100110011001,
0100110111111001100110011001,
0100111000001001100110011001,
0100111000011001100110011001,
0100111000101001100110011001,
0100111000111001100110011001,
0100111001001001100110011001,
0100111001011001100110011001,
0100111001101001100110011001,
0100111001111001100110011001,
0100111010001001100110011001,
0100111010011001100110011001,
0100111010101001100110011001,
0100111010111001100110011001,
0100111011001001100110011001,
0100111011011001100110011001,
0100111011101001100110011001,
0100111011111001100110011001,
0100111100001001100110011001,
0100111100011001100110011001,
0100111100101001100110011001,
0100111100111001100110011001,
0100111101001001100110011001,
0100111101011001100110011001,
0100111101101001100110011001,
0100111101111001100110011001,
0100111110001001100110011001,
0100111110011001100110011001,
0100111110101001100110011001,
0100111110111001100110011001,
0100111111001001100110011001,
0100111111011001100110011001,
0100111111101001100110011001,
0100111111111001100110011001,
0101000000001001100110011001,
0101000000011001100110011001,
0101000000101001100110011001,
0101000000111001100110011001,
0101000001001001100110011001,
0101000001011001100110011001,
0101000001101001100110011001,
0101000001111001100110011001,
0101000010001001100110011001,
0101000010011001100110011001,
0101000010101001100110011001,
0101000010111001100110011001,
0101000011001001100110011001,
0101000011011001100110011001,
0101000011101001100110011001,
0101000011111001100110011001,
0101000100001001100110011001,
0101000100011001100110011001,
0101000100101001100110011001,
0101000100111001100110011001,
0101000101001001100110011001,
0101000101011001100110011001,
0101000101101001100110011001,
0101000101111001100110011001,
0101000110001001100110011001,
0101000110011001100110011001,
0101000110101001100110011001,
0101000110111001100110011001,
0101000111001001100110011001,
0101000111011001100110011001,
0101000111101001100110011001,
0101000111111001100110011001,
0101001000001001100110011001,
0101001000011001100110011001,
0101001000101001100110011001,
0101001000111001100110011001,
0101001001001001100110011001,
0101001001011001100110011001,
0101001001101001100110011001,
0101001001111001100110011001,
0101001010001001100110011001,
0101001010011001100110011001,
0101001010101001100110011001,
0101001010111001100110011001,
0101001011001001100110011001,
0101001011011001100110011001,
0101001011101001100110011001,
0101001011111001100110011001,
0101001100001001100110011001,
0101001100011001100110011001,
0101001100101001100110011001,
0101001100111001100110011001,
0101001101001001100110011001,
0101001101011001100110011001,
0101001101101001100110011001,
0101001101111001100110011001,
0101001110001001100110011001,
0101001110011001100110011001,
0101001110101001100110011001,
0101001110111001100110011001,
0101001111001001100110011001,
0101001111011001100110011001,
0101001111101001100110011001,
0101001111111001100110011001,
0101010000001001100110011001,
0101010000011001100110011001,
0101010000101001100110011001,
0101010000111001100110011001,
0101010001001001100110011001,
0101010001011001100110011001,
0101010001101001100110011001,
0101010001111001100110011001,
0101010010001001100110011001,
0101010010011001100110011001,
0101010010101001100110011001,
0101010010111001100110011001,
0101010011001001100110011001,
0101010011011001100110011001,
0101010011101001100110011001,
0101010011111001100110011001,
0101010100001001100110011001,
0101010100011001100110011001,
0101010100101001100110011001,
0101010100111001100110011001,
0101010101001001100110011001,
0101010101011001100110011001,
0101010101101001100110011001,
0101010101111001100110011001,
0101010110001001100110011001,
0101010110011001100110011001,
0101010110101001100110011001,
0101010110111001100110011001,
0101010111001001100110011001,
0101010111011001100110011001,
0101010111101001100110011001,
0101010111111001100110011001,
0101011000001001100110011001,
0101011000011001100110011001,
0101011000101001100110011001,
0101011000111001100110011001,
0101011001001001100110011001,
0101011001011001100110011001,
0101011001101001100110011001,
0101011001111001100110011001,
0101011010001001100110011001,
0101011010011001100110011001,
0101011010101001100110011001,
0101011010111001100110011001,
0101011011001001100110011001,
0101011011011001100110011001,
0101011011101001100110011001,
0101011011111001100110011001,
0101011100001001100110011001,
0101011100011001100110011001,
0101011100101001100110011001,
0101011100111001100110011001,
0101011101001001100110011001,
0101011101011001100110011001,
0101011101101001100110011001,
0101011101111001100110011001,
0101011110001001100110011001,
0101011110011001100110011001,
0101011110101001100110011001,
0101011110111001100110011001,
0101011111001001100110011001,
0101011111011001100110011001,
0101011111101001100110011001,
0101011111111001100110011001,
0101100000001001100110011001,
0101100000011001100110011001,
0101100000101001100110011001,
0101100000111001100110011001,
0101100001001001100110011001,
0101100001011001100110011001,
0101100001101001100110011001,
0101100001111001100110011001,
0101100010001001100110011001,
0101100010011001100110011001,
0101100010101001100110011001,
0101100010111001100110011001,
0101100011001001100110011001,
0101100011011001100110011001,
0101100011101001100110011001,
0101100011111001100110011001,
0101100100001001100110011001,
0101100100011001100110011001,
0101100100101001100110011001,
0101100100111001100110011001,
0101100101001001100110011001,
0101100101011001100110011001,
0101100101101001100110011001,
0101100101111001100110011001,
0101100110001001100110011001,
0101100110011001100110011001,
0101100110101001100110011001,
0101100110111001100110011001,
0101100111001001100110011001,
0101100111011001100110011001,
0101100111101001100110011001,
0101100111111001100110011001,
0101101000001001100110011001,
0101101000011001100110011001,
0101101000101001100110011001,
0101101000111001100110011001,
0101101001001001100110011001,
0101101001011001100110011001,
0101101001101001100110011001,
0101101001111001100110011001,
0101101010001001100110011001,
0101101010011001100110011001,
0101101010101001100110011001,
0101101010111001100110011001,
0101101011001001100110011001,
0101101011011001100110011001,
0101101011101001100110011001,
0101101011111001100110011001,
0101101100001001100110011001,
0101101100011001100110011001,
0101101100101001100110011001,
0101101100111001100110011001,
0101101101001001100110011001,
0101101101011001100110011001,
0101101101101001100110011001,
0101101101111001100110011001,
0101101110001001100110011001,
0101101110011001100110011001,
0101101110101001100110011001,
0101101110111001100110011001,
0101101111001001100110011001,
0101101111011001100110011001,
0101101111101001100110011001,
0101101111111001100110011001,
0101110000001001100110011001,
0101110000011001100110011001,
0101110000101001100110011001,
0101110000111001100110011001,
0101110001001001100110011001,
0101110001011001100110011001,
0101110001101001100110011001,
0101110001111001100110011001,
0101110010001001100110011001,
0101110010011001100110011001,
0101110010101001100110011001,
0101110010111001100110011001,
0101110011001001100110011001,
0101110011011001100110011001,
0101110011101001100110011001,
0101110011111001100110011001,
0101110100001001100110011001,
0101110100011001100110011001,
0101110100101001100110011001,
0101110100111001100110011001,
0101110101001001100110011001,
0101110101011001100110011001,
0101110101101001100110011001,
0101110101111001100110011001,
0101110110001001100110011001,
0101110110011001100110011001,
0101110110101001100110011001,
0101110110111001100110011001,
0101110111001001100110011001,
0101110111011001100110011001,
0101110111101001100110011001,
0101110111111001100110011001,
0101111000001001100110011001,
0101111000011001100110011001,
0101111000101001100110011001,
0101111000111001100110011001,
0101111001001001100110011001,
0101111001011001100110011001,
0101111001101001100110011001,
0101111001111001100110011001,
0101111010001001100110011001,
0101111010011001100110011001,
0101111010101001100110011001,
0101111010111001100110011001,
0101111011001001100110011001,
0101111011011001100110011001,
0101111011101001100110011001,
0101111011111001100110011001,
0101111100001001100110011001,
0101111100011001100110011001,
0101111100101001100110011001,
0101111100111001100110011001,
0101111101001001100110011001,
0101111101011001100110011001,
0101111101101001100110011001,
0101111101111001100110011001,
0101111110001001100110011001,
0101111110011001100110011001,
0101111110101001100110011001,
0101111110111001100110011001,
0101111111001001100110011001,
0101111111011001100110011001,
0101111111101001100110011001,
0101111111111001100110011001,
0110000000001001100110011001,
0110000000011001100110011001,
0110000000101001100110011001,
0110000000111001100110011001,
0110000001001001100110011001,
0110000001011001100110011001,
0110000001101001100110011001,
0110000001111001100110011001,
0110000010001001100110011001,
0110000010011001100110011001,
0110000010101001100110011001,
0110000010111001100110011001,
0110000011001001100110011001,
0110000011011001100110011001,
0110000011101001100110011001,
0110000011111001100110011001,
0110000100001001100110011001,
0110000100011001100110011001,
0110000100101001100110011001,
0110000100111001100110011001,
0110000101001001100110011001,
0110000101011001100110011001,
0110000101101001100110011001,
0110000101111001100110011001,
0110000110001001100110011001,
0110000110011001100110011001,
0110000110101001100110011001,
0110000110111001100110011001,
0110000111001001100110011001,
0110000111011001100110011001,
0110000111101001100110011001,
0110000111111001100110011001,
0110001000001001100110011001,
0110001000011001100110011001,
0110001000101001100110011001,
0110001000111001100110011001,
0110001001001001100110011001,
0110001001011001100110011001,
0110001001101001100110011001,
0110001001111001100110011001,
0110001010001001100110011001,
0110001010011001100110011001,
0110001010101001100110011001,
0110001010111001100110011001,
0110001011001001100110011001,
0110001011011001100110011001,
0110001011101001100110011001,
0110001011111001100110011001,
0110001100001001100110011001,
0110001100011001100110011001,
0110001100101001100110011001,
0110001100111001100110011001,
0110001101001001100110011001,
0110001101011001100110011001,
0110001101101001100110011001,
0110001101111001100110011001,
0110001110001001100110011001,
0110001110011001100110011001,
0110001110101001100110011001,
0110001110111001100110011001,
0110001111001001100110011001,
0110001111011001100110011001,
0110001111101001100110011001,
0110001111111001100110011001,
0110010000001001100110011001,
0110010000011001100110011001,
0110010000101001100110011001,
0110010000111001100110011001,
0110010001001001100110011001,
0110010001011001100110011001,
0110010001101001100110011001,
0110010001111001100110011001,
0110010010001001100110011001,
0110010010011001100110011001,
0110010010101001100110011001,
0110010010111001100110011001,
0110010011001001100110011001,
0110010011011001100110011001,
0110010011101001100110011001,
0110010011111001100110011001,
0110010100001001100110011001,
0110010100011001100110011001,
0110010100101001100110011001,
0110010100111001100110011001,
0110010101001001100110011001,
0110010101011001100110011001,
0110010101101001100110011001,
0110010101111001100110011001,
0110010110001001100110011001,
0110010110011001100110011001,
0110010110101001100110011001,
0110010110111001100110011001,
0110010111001001100110011001,
0110010111011001100110011001,
0110010111101001100110011001,
0110010111111001100110011001,
0110011000001001100110011001,
0110011000011001100110011001,
0110011000101001100110011001,
0110011000111001100110011001,
0110011001001001100110011001,
0110011001011001100110011001,
0110011001101001100110011001,
0110011001111001100110011001,
0110011010001001100110011001,
0110011010011001100110011001,
0110011010101001100110011001,
0110011010111001100110011001,
0110011011001001100110011001,
0110011011011001100110011001,
0110011011101001100110011001,
0110011011111001100110011001,
0110011100001001100110011001,
0110011100011001100110011001,
0110011100101001100110011001,
0110011100111001100110011001,
0110011101001001100110011001,
0110011101011001100110011001,
0110011101101001100110011001,
0110011101111001100110011001,
0110011110001001100110011001,
0110011110011001100110011001,
0110011110101001100110011001,
0110011110111001100110011001,
0110011111001001100110011001,
0110011111011001100110011001,
0110011111101001100110011001,
0110011111111001100110011001,
0110100000001001100110011001,
0110100000011001100110011001,
0110100000101001100110011001,
0110100000111001100110011001,
0110100001001001100110011001,
0110100001011001100110011001,
0110100001101001100110011001,
0110100001111001100110011001,
0110100010001001100110011001,
0110100010011001100110011001,
0110100010101001100110011001,
0110100010111001100110011001,
0110100011001001100110011001,
0110100011011001100110011001,
0110100011101001100110011001,
0110100011111001100110011001,
0110100100001001100110011001,
0110100100011001100110011001,
0110100100101001100110011001,
0110100100111001100110011001,
0110100101001001100110011001,
0110100101011001100110011001,
0110100101101001100110011001,
0110100101111001100110011001,
0110100110001001100110011001,
0110100110011001100110011001,
0110100110101001100110011001,
0110100110111001100110011001,
0110100111001001100110011001,
0110100111011001100110011001,
0110100111101001100110011001,
0110100111111001100110011001,
0110101000001001100110011001,
0110101000011001100110011001,
0110101000101001100110011001,
0110101000111001100110011001,
0110101001001001100110011001,
0110101001011001100110011001,
0110101001101001100110011001,
0110101001111001100110011001,
0110101010001001100110011001,
0110101010011001100110011001,
0110101010101001100110011001,
0110101010111001100110011001,
0110101011001001100110011001,
0110101011011001100110011001,
0110101011101001100110011001,
0110101011111001100110011001,
0110101100001001100110011001,
0110101100011001100110011001,
0110101100101001100110011001,
0110101100111001100110011001,
0110101101001001100110011001,
0110101101011001100110011001,
0110101101101001100110011001,
0110101101111001100110011001,
0110101110001001100110011001,
0110101110011001100110011001,
0110101110101001100110011001,
0110101110111001100110011001,
0110101111001001100110011001,
0110101111011001100110011001,
0110101111101001100110011001,
0110101111111001100110011001,
0110110000001001100110011001,
0110110000011001100110011001,
0110110000101001100110011001,
0110110000111001100110011001,
0110110001001001100110011001,
0110110001011001100110011001,
0110110001101001100110011001,
0110110001111001100110011001,
0110110010001001100110011001,
0110110010011001100110011001,
0110110010101001100110011001,
0110110010111001100110011001,
0110110011001001100110011001,
0110110011011001100110011001,
0110110011101001100110011001,
0110110011111001100110011001,
0110110100001001100110011001,
0110110100011001100110011001,
0110110100101001100110011001,
0110110100111001100110011001,
0110110101001001100110011001,
0110110101011001100110011001,
0110110101101001100110011001,
0110110101111001100110011001,
0110110110001001100110011001,
0110110110011001100110011001,
0110110110101001100110011001,
0110110110111001100110011001,
0110110111001001100110011001,
0110110111011001100110011001,
0110110111101001100110011001,
0110110111111001100110011001,
0110111000001001100110011001,
0110111000011001100110011001,
0110111000101001100110011001,
0110111000111001100110011001,
0110111001001001100110011001,
0110111001011001100110011001,
0110111001101001100110011001,
0110111001111001100110011001,
0110111010001001100110011001,
0110111010011001100110011001,
0110111010101001100110011001,
0110111010111001100110011001,
0110111011001001100110011001,
0110111011011001100110011001,
0110111011101001100110011001,
0110111011111001100110011001,
0110111100001001100110011001,
0110111100011001100110011001,
0110111100101001100110011001,
0110111100111001100110011001,
0110111101001001100110011001,
0110111101011001100110011001,
0110111101101001100110011001,
0110111101111001100110011001,
0110111110001001100110011001,
0110111110011001100110011001,
0110111110101001100110011001,
0110111110111001100110011001,
0110111111001001100110011001,
0110111111011001100110011001,
0110111111101001100110011001,
0110111111111001100110011001,
0111000000001001100110011001,
0111000000011001100110011001,
0111000000101001100110011001,
0111000000111001100110011001,
0111000001001001100110011001,
0111000001011001100110011001,
0111000001101001100110011001,
0111000001111001100110011001,
0111000010001001100110011001,
0111000010011001100110011001,
0111000010101001100110011001,
0111000010111001100110011001,
0111000011001001100110011001,
0111000011011001100110011001,
0111000011101001100110011001,
0111000011111001100110011001,
0111000100001001100110011001,
0111000100011001100110011001,
0111000100101001100110011001,
0111000100111001100110011001,
0111000101001001100110011001,
0111000101011001100110011001,
0111000101101001100110011001,
0111000101111001100110011001,
0111000110001001100110011001,
0111000110011001100110011001,
0111000110101001100110011001,
0111000110111001100110011001,
0111000111001001100110011001,
0111000111011001100110011001,
0111000111101001100110011001,
0111000111111001100110011001,
0111001000001001100110011001,
0111001000011001100110011001,
0111001000101001100110011001,
0111001000111001100110011001,
0111001001001001100110011001,
0111001001011001100110011001,
0111001001101001100110011001,
0111001001111001100110011001,
0111001010001001100110011001,
0111001010011001100110011001,
0111001010101001100110011001,
0111001010111001100110011001,
0111001011001001100110011001,
0111001011011001100110011001,
0111001011101001100110011001,
0111001011111001100110011001,
0111001100001001100110011001,
0111001100011001100110011001,
0111001100101001100110011001,
0111001100111001100110011001,
0111001101001001100110011001,
0111001101011001100110011001,
0111001101101001100110011001,
0111001101111001100110011001,
0111001110001001100110011001,
0111001110011001100110011001,
0111001110101001100110011001,
0111001110111001100110011001,
0111001111001001100110011001,
0111001111011001100110011001,
0111001111101001100110011001,
0111001111111001100110011001,
0111010000001001100110011001,
0111010000011001100110011001,
0111010000101001100110011001,
0111010000111001100110011001,
0111010001001001100110011001,
0111010001011001100110011001,
0111010001101001100110011001,
0111010001111001100110011001,
0111010010001001100110011001,
0111010010011001100110011001,
0111010010101001100110011001,
0111010010111001100110011001,
0111010011001001100110011001,
0111010011011001100110011001,
0111010011101001100110011001,
0111010011111001100110011001,
0111010100001001100110011001,
0111010100011001100110011001,
0111010100101001100110011001,
0111010100111001100110011001,
0111010101001001100110011001,
0111010101011001100110011001,
0111010101101001100110011001,
0111010101111001100110011001,
0111010110001001100110011001,
0111010110011001100110011001,
0111010110101001100110011001,
0111010110111001100110011001,
0111010111001001100110011001,
0111010111011001100110011001,
0111010111101001100110011001,
0111010111111001100110011001,
0111011000001001100110011001,
0111011000011001100110011001,
0111011000101001100110011001,
0111011000111001100110011001,
0111011001001001100110011001,
0111011001011001100110011001,
0111011001101001100110011001,
0111011001111001100110011001,
0111011010001001100110011001,
0111011010011001100110011001,
0111011010101001100110011001,
0111011010111001100110011001,
0111011011001001100110011001,
0111011011011001100110011001,
0111011011101001100110011001,
0111011011111001100110011001,
0111011100001001100110011001,
0111011100011001100110011001,
0111011100101001100110011001,
0111011100111001100110011001,
0111011101001001100110011001,
0111011101011001100110011001,
0111011101101001100110011001,
0111011101111001100110011001,
0111011110001001100110011001,
0111011110011001100110011001,
0111011110101001100110011001,
0111011110111001100110011001,
0111011111001001100110011001,
0111011111011001100110011001,
0111011111101001100110011001,
0111011111111001100110011001,
0111100000001001100110011001,
0111100000011001100110011001,
0111100000101001100110011001,
0111100000111001100110011001,
0111100001001001100110011001,
0111100001011001100110011001,
0111100001101001100110011001,
0111100001111001100110011001,
0111100010001001100110011001,
0111100010011001100110011001,
0111100010101001100110011001,
0111100010111001100110011001,
0111100011001001100110011001,
0111100011011001100110011001,
0111100011101001100110011001,
0111100011111001100110011001,
0111100100001001100110011001,
0111100100011001100110011001,
0111100100101001100110011001,
0111100100111001100110011001,
0111100101001001100110011001,
0111100101011001100110011001,
0111100101101001100110011001,
0111100101111001100110011001,
0111100110001001100110011001,
0111100110011001100110011001,
0111100110101001100110011001,
0111100110111001100110011001,
0111100111001001100110011001,
0111100111011001100110011001,
0111100111101001100110011001,
0111100111111001100110011001,
0111101000001001100110011001,
0111101000011001100110011001,
0111101000101001100110011001,
0111101000111001100110011001,
0111101001001001100110011001,
0111101001011001100110011001,
0111101001101001100110011001,
0111101001111001100110011001,
0111101010001001100110011001,
0111101010011001100110011001,
0111101010101001100110011001,
0111101010111001100110011001,
0111101011001001100110011001,
0111101011011001100110011001,
0111101011101001100110011001,
0111101011111001100110011001,
0111101100001001100110011001,
0111101100011001100110011001,
0111101100101001100110011001,
0111101100111001100110011001,
0111101101001001100110011001,
0111101101011001100110011001,
0111101101101001100110011001,
0111101101111001100110011001,
0111101110001001100110011001,
0111101110011001100110011001,
0111101110101001100110011001,
0111101110111001100110011001,
0111101111001001100110011001,
0111101111011001100110011001,
0111101111101001100110011001,
0111101111111001100110011001,
0111110000001001100110011001,
0111110000011001100110011001,
0111110000101001100110011001,
0111110000111001100110011001,
0111110001001001100110011001,
0111110001011001100110011001,
0111110001101001100110011001,
0111110001111001100110011001,
0111110010001001100110011001,
0111110010011001100110011001,
0111110010101001100110011001,
0111110010111001100110011001,
0111110011001001100110011001,
0111110011011001100110011001,
0111110011101001100110011001,
0111110011111001100110011001,
0111110100001001100110011001,
0111110100011001100110011001,
0111110100101001100110011001,
0111110100111001100110011001,
0111110101001001100110011001,
0111110101011001100110011001,
0111110101101001100110011001,
0111110101111001100110011001,
0111110110001001100110011001,
0111110110011001100110011001,
0111110110101001100110011001,
0111110110111001100110011001,
0111110111001001100110011001,
0111110111011001100110011001,
0111110111101001100110011001,
0111110111111001100110011001,
0111111000001001100110011001,
0111111000011001100110011001,
0111111000101001100110011001,
0111111000111001100110011001,
0111111001001001100110011001,
0111111001011001100110011001,
0111111001101001100110011001,
0111111001111001100110011001,
0111111010001001100110011001,
0111111010011001100110011001,
0111111010101001100110011001,
0111111010111001100110011001,
0111111011001001100110011001,
0111111011011001100110011001,
0111111011101001100110011001,
0111111011111001100110011001,
0111111100001001100110011001,
0111111100011001100110011001,
0111111100101001100110011001,
0111111100111001100110011001,
0111111101001001100110011001,
0111111101011001100110011001,
0111111101101001100110011001,
0111111101111001100110011001,
0111111110001001100110011001,
0111111110011001100110011001,
0111111110101001100110011001,
0111111110111001100110011001,
0111111111001001100110011001,
0111111111011001100110011001,
0111111111101001100110011001,
0111111111111001100110011001
);

type muon_pt_lut_array is array (0 to 2**(D_S_I_MUON_V2.pt_high-D_S_I_MUON_V2.pt_low+1)-1) of sfixed(9 downto -17);

constant MU_PT_LUT_SFIXED : muon_pt_lut_array := (
00000000000000000000000000,
00000000001001100110011001,
00000000011001100110011001,
00000000101001100110011001,
00000000111001100110011001,
00000001001001100110011001,
00000001011001100110011001,
00000001101001100110011001,
00000001111001100110011001,
00000010001001100110011001,
00000010011001100110011001,
00000010101001100110011001,
00000010111001100110011001,
00000011001001100110011001,
00000011011001100110011001,
00000011101001100110011001,
00000011111001100110011001,
00000100001001100110011001,
00000100011001100110011001,
00000100101001100110011001,
00000100111001100110011001,
00000101001001100110011001,
00000101011001100110011001,
00000101101001100110011001,
00000101111001100110011001,
00000110001001100110011001,
00000110011001100110011001,
00000110101001100110011001,
00000110111001100110011001,
00000111001001100110011001,
00000111011001100110011001,
00000111101001100110011001,
00000111111001100110011001,
00001000001001100110011001,
00001000011001100110011001,
00001000101001100110011001,
00001000111001100110011001,
00001001001001100110011001,
00001001011001100110011001,
00001001101001100110011001,
00001001111001100110011001,
00001010001001100110011001,
00001010011001100110011001,
00001010101001100110011001,
00001010111001100110011001,
00001011001001100110011001,
00001011011001100110011001,
00001011101001100110011001,
00001011111001100110011001,
00001100001001100110011001,
00001100011001100110011001,
00001100101001100110011001,
00001100111001100110011001,
00001101001001100110011001,
00001101011001100110011001,
00001101101001100110011001,
00001101111001100110011001,
00001110001001100110011001,
00001110011001100110011001,
00001110101001100110011001,
00001110111001100110011001,
00001111001001100110011001,
00001111011001100110011001,
00001111101001100110011001,
00001111111001100110011001,
00010000001001100110011001,
00010000011001100110011001,
00010000101001100110011001,
00010000111001100110011001,
00010001001001100110011001,
00010001011001100110011001,
00010001101001100110011001,
00010001111001100110011001,
00010010001001100110011001,
00010010011001100110011001,
00010010101001100110011001,
00010010111001100110011001,
00010011001001100110011001,
00010011011001100110011001,
00010011101001100110011001,
00010011111001100110011001,
00010100001001100110011001,
00010100011001100110011001,
00010100101001100110011001,
00010100111001100110011001,
00010101001001100110011001,
00010101011001100110011001,
00010101101001100110011001,
00010101111001100110011001,
00010110001001100110011001,
00010110011001100110011001,
00010110101001100110011001,
00010110111001100110011001,
00010111001001100110011001,
00010111011001100110011001,
00010111101001100110011001,
00010111111001100110011001,
00011000001001100110011001,
00011000011001100110011001,
00011000101001100110011001,
00011000111001100110011001,
00011001001001100110011001,
00011001011001100110011001,
00011001101001100110011001,
00011001111001100110011001,
00011010001001100110011001,
00011010011001100110011001,
00011010101001100110011001,
00011010111001100110011001,
00011011001001100110011001,
00011011011001100110011001,
00011011101001100110011001,
00011011111001100110011001,
00011100001001100110011001,
00011100011001100110011001,
00011100101001100110011001,
00011100111001100110011001,
00011101001001100110011001,
00011101011001100110011001,
00011101101001100110011001,
00011101111001100110011001,
00011110001001100110011001,
00011110011001100110011001,
00011110101001100110011001,
00011110111001100110011001,
00011111001001100110011001,
00011111011001100110011001,
00011111101001100110011001,
00011111111001100110011001,
00100000001001100110011001,
00100000011001100110011001,
00100000101001100110011001,
00100000111001100110011001,
00100001001001100110011001,
00100001011001100110011001,
00100001101001100110011001,
00100001111001100110011001,
00100010001001100110011001,
00100010011001100110011001,
00100010101001100110011001,
00100010111001100110011001,
00100011001001100110011001,
00100011011001100110011001,
00100011101001100110011001,
00100011111001100110011001,
00100100001001100110011001,
00100100011001100110011001,
00100100101001100110011001,
00100100111001100110011001,
00100101001001100110011001,
00100101011001100110011001,
00100101101001100110011001,
00100101111001100110011001,
00100110001001100110011001,
00100110011001100110011001,
00100110101001100110011001,
00100110111001100110011001,
00100111001001100110011001,
00100111011001100110011001,
00100111101001100110011001,
00100111111001100110011001,
00101000001001100110011001,
00101000011001100110011001,
00101000101001100110011001,
00101000111001100110011001,
00101001001001100110011001,
00101001011001100110011001,
00101001101001100110011001,
00101001111001100110011001,
00101010001001100110011001,
00101010011001100110011001,
00101010101001100110011001,
00101010111001100110011001,
00101011001001100110011001,
00101011011001100110011001,
00101011101001100110011001,
00101011111001100110011001,
00101100001001100110011001,
00101100011001100110011001,
00101100101001100110011001,
00101100111001100110011001,
00101101001001100110011001,
00101101011001100110011001,
00101101101001100110011001,
00101101111001100110011001,
00101110001001100110011001,
00101110011001100110011001,
00101110101001100110011001,
00101110111001100110011001,
00101111001001100110011001,
00101111011001100110011001,
00101111101001100110011001,
00101111111001100110011001,
00110000001001100110011001,
00110000011001100110011001,
00110000101001100110011001,
00110000111001100110011001,
00110001001001100110011001,
00110001011001100110011001,
00110001101001100110011001,
00110001111001100110011001,
00110010001001100110011001,
00110010011001100110011001,
00110010101001100110011001,
00110010111001100110011001,
00110011001001100110011001,
00110011011001100110011001,
00110011101001100110011001,
00110011111001100110011001,
00110100001001100110011001,
00110100011001100110011001,
00110100101001100110011001,
00110100111001100110011001,
00110101001001100110011001,
00110101011001100110011001,
00110101101001100110011001,
00110101111001100110011001,
00110110001001100110011001,
00110110011001100110011001,
00110110101001100110011001,
00110110111001100110011001,
00110111001001100110011001,
00110111011001100110011001,
00110111101001100110011001,
00110111111001100110011001,
00111000001001100110011001,
00111000011001100110011001,
00111000101001100110011001,
00111000111001100110011001,
00111001001001100110011001,
00111001011001100110011001,
00111001101001100110011001,
00111001111001100110011001,
00111010001001100110011001,
00111010011001100110011001,
00111010101001100110011001,
00111010111001100110011001,
00111011001001100110011001,
00111011011001100110011001,
00111011101001100110011001,
00111011111001100110011001,
00111100001001100110011001,
00111100011001100110011001,
00111100101001100110011001,
00111100111001100110011001,
00111101001001100110011001,
00111101011001100110011001,
00111101101001100110011001,
00111101111001100110011001,
00111110001001100110011001,
00111110011001100110011001,
00111110101001100110011001,
00111110111001100110011001,
00111111001001100110011001,
00111111011001100110011001,
00111111101001100110011001,
00111111111001100110011001,
01000000001001100110011001,
01000000011001100110011001,
01000000101001100110011001,
01000000111001100110011001,
01000001001001100110011001,
01000001011001100110011001,
01000001101001100110011001,
01000001111001100110011001,
01000010001001100110011001,
01000010011001100110011001,
01000010101001100110011001,
01000010111001100110011001,
01000011001001100110011001,
01000011011001100110011001,
01000011101001100110011001,
01000011111001100110011001,
01000100001001100110011001,
01000100011001100110011001,
01000100101001100110011001,
01000100111001100110011001,
01000101001001100110011001,
01000101011001100110011001,
01000101101001100110011001,
01000101111001100110011001,
01000110001001100110011001,
01000110011001100110011001,
01000110101001100110011001,
01000110111001100110011001,
01000111001001100110011001,
01000111011001100110011001,
01000111101001100110011001,
01000111111001100110011001,
01001000001001100110011001,
01001000011001100110011001,
01001000101001100110011001,
01001000111001100110011001,
01001001001001100110011001,
01001001011001100110011001,
01001001101001100110011001,
01001001111001100110011001,
01001010001001100110011001,
01001010011001100110011001,
01001010101001100110011001,
01001010111001100110011001,
01001011001001100110011001,
01001011011001100110011001,
01001011101001100110011001,
01001011111001100110011001,
01001100001001100110011001,
01001100011001100110011001,
01001100101001100110011001,
01001100111001100110011001,
01001101001001100110011001,
01001101011001100110011001,
01001101101001100110011001,
01001101111001100110011001,
01001110001001100110011001,
01001110011001100110011001,
01001110101001100110011001,
01001110111001100110011001,
01001111001001100110011001,
01001111011001100110011001,
01001111101001100110011001,
01001111111001100110011001,
01010000001001100110011001,
01010000011001100110011001,
01010000101001100110011001,
01010000111001100110011001,
01010001001001100110011001,
01010001011001100110011001,
01010001101001100110011001,
01010001111001100110011001,
01010010001001100110011001,
01010010011001100110011001,
01010010101001100110011001,
01010010111001100110011001,
01010011001001100110011001,
01010011011001100110011001,
01010011101001100110011001,
01010011111001100110011001,
01010100001001100110011001,
01010100011001100110011001,
01010100101001100110011001,
01010100111001100110011001,
01010101001001100110011001,
01010101011001100110011001,
01010101101001100110011001,
01010101111001100110011001,
01010110001001100110011001,
01010110011001100110011001,
01010110101001100110011001,
01010110111001100110011001,
01010111001001100110011001,
01010111011001100110011001,
01010111101001100110011001,
01010111111001100110011001,
01011000001001100110011001,
01011000011001100110011001,
01011000101001100110011001,
01011000111001100110011001,
01011001001001100110011001,
01011001011001100110011001,
01011001101001100110011001,
01011001111001100110011001,
01011010001001100110011001,
01011010011001100110011001,
01011010101001100110011001,
01011010111001100110011001,
01011011001001100110011001,
01011011011001100110011001,
01011011101001100110011001,
01011011111001100110011001,
01011100001001100110011001,
01011100011001100110011001,
01011100101001100110011001,
01011100111001100110011001,
01011101001001100110011001,
01011101011001100110011001,
01011101101001100110011001,
01011101111001100110011001,
01011110001001100110011001,
01011110011001100110011001,
01011110101001100110011001,
01011110111001100110011001,
01011111001001100110011001,
01011111011001100110011001,
01011111101001100110011001,
01011111111001100110011001,
01100000001001100110011001,
01100000011001100110011001,
01100000101001100110011001,
01100000111001100110011001,
01100001001001100110011001,
01100001011001100110011001,
01100001101001100110011001,
01100001111001100110011001,
01100010001001100110011001,
01100010011001100110011001,
01100010101001100110011001,
01100010111001100110011001,
01100011001001100110011001,
01100011011001100110011001,
01100011101001100110011001,
01100011111001100110011001,
01100100001001100110011001,
01100100011001100110011001,
01100100101001100110011001,
01100100111001100110011001,
01100101001001100110011001,
01100101011001100110011001,
01100101101001100110011001,
01100101111001100110011001,
01100110001001100110011001,
01100110011001100110011001,
01100110101001100110011001,
01100110111001100110011001,
01100111001001100110011001,
01100111011001100110011001,
01100111101001100110011001,
01100111111001100110011001,
01101000001001100110011001,
01101000011001100110011001,
01101000101001100110011001,
01101000111001100110011001,
01101001001001100110011001,
01101001011001100110011001,
01101001101001100110011001,
01101001111001100110011001,
01101010001001100110011001,
01101010011001100110011001,
01101010101001100110011001,
01101010111001100110011001,
01101011001001100110011001,
01101011011001100110011001,
01101011101001100110011001,
01101011111001100110011001,
01101100001001100110011001,
01101100011001100110011001,
01101100101001100110011001,
01101100111001100110011001,
01101101001001100110011001,
01101101011001100110011001,
01101101101001100110011001,
01101101111001100110011001,
01101110001001100110011001,
01101110011001100110011001,
01101110101001100110011001,
01101110111001100110011001,
01101111001001100110011001,
01101111011001100110011001,
01101111101001100110011001,
01101111111001100110011001,
01110000001001100110011001,
01110000011001100110011001,
01110000101001100110011001,
01110000111001100110011001,
01110001001001100110011001,
01110001011001100110011001,
01110001101001100110011001,
01110001111001100110011001,
01110010001001100110011001,
01110010011001100110011001,
01110010101001100110011001,
01110010111001100110011001,
01110011001001100110011001,
01110011011001100110011001,
01110011101001100110011001,
01110011111001100110011001,
01110100001001100110011001,
01110100011001100110011001,
01110100101001100110011001,
01110100111001100110011001,
01110101001001100110011001,
01110101011001100110011001,
01110101101001100110011001,
01110101111001100110011001,
01110110001001100110011001,
01110110011001100110011001,
01110110101001100110011001,
01110110111001100110011001,
01110111001001100110011001,
01110111011001100110011001,
01110111101001100110011001,
01110111111001100110011001,
01111000001001100110011001,
01111000011001100110011001,
01111000101001100110011001,
01111000111001100110011001,
01111001001001100110011001,
01111001011001100110011001,
01111001101001100110011001,
01111001111001100110011001,
01111010001001100110011001,
01111010011001100110011001,
01111010101001100110011001,
01111010111001100110011001,
01111011001001100110011001,
01111011011001100110011001,
01111011101001100110011001,
01111011111001100110011001,
01111100001001100110011001,
01111100011001100110011001,
01111100101001100110011001,
01111100111001100110011001,
01111101001001100110011001,
01111101011001100110011001,
01111101101001100110011001,
01111101111001100110011001,
01111110001001100110011001,
01111110011001100110011001,
01111110101001100110011001,
01111110111001100110011001,
01111111001001100110011001,
01111111011001100110011001,
01111111101001100110011001
);

-- calo-calo cosh deta LUTs
type calo_calo_cosh_deta_lut_sfixed_array is array (0 to 2**MAX_CALO_ETA_BITS-1) of sfixed(15 downto -19);

constant CALO_CALO_COSH_DETA_LUT_SFIXED : calo_calo_cosh_deta_lut_sfixed_array := (
0000000000000010000000000000000000,
0000000000000010000000001000001100,
0000000000000010000000100000110001,
0000000000000010000001001001101110,
0000000000000010000001111010111000,
0000000000000010000011000100100110,
0000000000000010000100010110100001,
0000000000000010000110000001000001,
0000000000000010000111110011101101,
0000000000000010001001111110111110,
0000000000000010001100010010011011,
0000000000000010001110111110011101,
0000000000000010010001110010101100,
0000000000000010010100111111011111,
0000000000000010011000011100101011,
0000000000000010011100010010011011,
0000000000000010100000010000011000,
0000000000000010100100100110111010,
0000000000000010101001010110000001,
0000000000000010101110001101010011,
0000000000000010110011100101011000,
0000000000000010111001001101110100,
0000000000000010111111001110110110,
0000000000000011000101101000011100,
0000000000000011001100010010011011,
0000000000000011010011011101001011,
0000000000000011011011000000100000,
0000000000000011100010111100011010,
0000000000000011101011010000111001,
0000000000000011110100000110001001,
0000000000000011111101010011111101,
0000000000000100000111001010110000,
0000000000000100010001011010000111,
0000000000000100011100001010001111,
0000000000000100100111011011001000,
0000000000000100110011010100111111,
0000000000000100111111101111100111,
0000000000000101001100110011001100,
0000000000000101011010011111101111,
0000000000000101101000110101001111,
0000000000000101110111110011101101,
0000000000000110000111100011010100,
0000000000000110011000000100000110,
0000000000000110101001010110000001,
0000000000000110111011011001000101,
0000000000000111001110001101010011,
0000000000000111100010000011000100,
0000000000000111110110101001111110,
0000000000001000001100010010011011,
0000000000001000100010111100011010,
0000000000001000111010100111111011,
0000000000001001010011010100111111,
0000000000001001101101001011110001,
0000000000001010001000001100010010,
0000000000001010100100011110101110,
0000000000001011000010000011000100,
0000000000001011100000111001010110,
0000000000001100000001010001111010,
0000000000001100100010111100011010,
0000000000001101000110001001001101,
0000000000001101101011000000100000,
0000000000001110010001100010010011,
0000000000001110111001101110100101,
0000000000001111100011110101110000,
0000000000010000001111101111100111,
0000000000010000111101100100010110,
0000000000010001101101100100010110,
0000000000010010011111100111011011,
0000000000010011010011111101111100,
0000000000010100001010100111111011,
0000000000010101000011101101100100,
0000000000010101111111010111000010,
0000000000010110111101101100100010,
0000000000010111111110101110000101,
0000000000011001000010110100001110,
0000000000011010001001110110110010,
0000000000011011010011111101111100,
0000000000011100100001100010010011,
0000000000011101110010011011101001,
0000000000011111000111000010100011,
0000000000100000011111010111000010,
0000000000100001111011101001011110,
0000000000100011011100000010000011,
0000000000100101000000110001001001,
0000000000100110101001110110110010,
0000000000101000010111110011101101,
0000000000101010001010011111101111,
0000000000101100000010010011011101,
0000000000101101111111011111001110,
0000000000110000000010010011011101,
0000000000110010001010111000010100,
0000000000110100011001011110001101,
0000000000110110101110011101101100,
0000000000111001001010000111001010,
0000000000111011101100100010110100,
0000000000111110010110011001100110,
0000000001000001000111101011100001,
0000000001000100000000111001010110,
0000000001000111000010010011011101,
0000000001001010001100011010100111,
0000000001001101011111011111001110,
0000000001010000111011111001110110,
0000000001010100100010000011000100,
0000000001011000010010100011110101,
0000000001011100001101101100100010,
0000000001100000010100000110001001,
0000000001100100100110000001000001,
0000000001101001000100001110010101,
0000000001101101101111000110101001,
0000000001110010100111010010111100,
0000000001110111101101011100001010,
0000000001111101000010000011000100,
0000000010000010100101110000101000,
0000000010001000011001001101110100,
0000000010001110011101010011111101,
0000000010010100110010101100000010,
0000000010011011011001111110111110,
0000000010100010010100000110001001,
0000000010101001100001111010111000,
0000000010110001000100010110100001,
0000000010111000111100001010001111,
0000000011000001001010010111100011,
0000000011001001101111111111111111,
0000000011010010101101111100111011,
0000000011011100000101100000010000,
0000000011100101110111110011101101,
0000000011110000000101110000101000,
0000000011111010110000111001010110,
0000000100000101111010011111101111,
0000000100010001100011101101100100,
0000000100011101101110000101000111,
0000000100101010011011000000100000,
0000000100110111101100001010001111,
0000000101000101100011000100100110,
0000000101010100000001011010000111,
0000000101100011001000110101001111,
0000000101110010111011011001000101,
0000000110000011011010110000001000,
0000000110010100101001001101110100,
0000000110100110101000100100110111,
0000000110111001011011001000101101,
0000000111001101000011001100110011,
0000000111100001100011000100100110,
0000000111110110111101001011110001,
0000001000001101010100010110100001,
0000001000100100101011001000101101,
0000001000111101000100010110100001,
0000001001010110100010111100011010,
0000001001110001001001111110111110,
0000001010001100111100111011011001,
0000001010101001111110110110010001,
0000001011001000010011010100111111,
0000001011100111111110000101000111,
0000001100001001000011000100100110,
0000001100101011100110001001001101,
0000001101001111101011011001000101,
0000001101110101010111011011001000,
0000001110011100101110101110000101,
0000001111000101110101111000110101,
0000001111110000110010001011010000,
0000010000011101101000100100110111,
0000010001001100011110101110000101,
0000010001111101011001111110111110,
0000010010110000100000100000110001,
0000010011100101111000100100110111,
0000010100011101101000010100011110,
0000010101010111110110110010001011,
0000010110010100101011000000100000,
0000010111010100001100001010001111,
0000011000010110100010001011010000,
0000011001011011110100110111010010,
0000011010100100001100101011000000,
0000011011101111110010100011110101,
0000011100111110101111010111000010,
0000011110010001001100111011011001,
0000011111100111010101000111101011,
0000100001000001010010011011101001,
0000100010011111001111100111011011,
0000100100000001011000001100010010,
0000100101100111111000000100000110,
0000100111010010111011100001010001,
0000101001000010101111100111011011,
0000101010110111100001110010101100,
0000101100110001100000011000100100,
0000101110110000111001111110111110,
0000110000110101111110000101000111,
0000110011000000111100111011011001,
0000110101010010000111000010100011,
0000110111101001101110010101100000,
0000111010001000000100111111011111,
0000111100101101011110010101100000,
0000111111011010001110001101010011,
0001000010001110101001100110011001,
0001000101001011000110011001100110,
0001001000001111111011011001000101,
0001001011011101100000100000110001,
0001001110110100001110100101111000,
0001010010010100011111101111100111,
0001010101111110101110110110010001,
0001011001110011011000100100110111,
0001011101110010111010010111100011,
0001100001111101110011010100111111,
0001100110010100100011101101100100,
0001101010110111101101001011110001,
0001101111100111110011001100110011,
0001110100100101011010010111100011,
0001111001110001001001010110000001,
0001111111001011101000010100011110,
0010000100110101100001001001101110,
0010001010101111011111101111100111,
0010010000111010010001110010101100,
0010010111010110100111001010110000,
0010011110000101010001110010101100,
0010100101000111000101111000110101,
0010101100011100111001111110111110,
0010110100000111100110110010001011,
0010111100001000000111111011111001,
0011000100011111011011011001000101,
0011001101001110100010000011000100,
0011010110010110011111011111001110,
0011011111111000011010100111111011,
0011101001110101011101010011111101,
0011110100001110110100100110111010,
0011111111000101110001001001101110,
0100001010011011100111001010110000,
0100010110010001101110011101101100,
0100100010101001100010111100011010,
0100101111100100100100100110111010,
0100111101000100010111011011001000,
0101001011001010100100000110001001,
0000000000000000000000000000000000,
0000000000000000000000000000000000,
0000000000000000000000000000000000,
0000000000000000000000000000000000,
0000000000000000000000000000000000,
0000000000000000000000000000000000,
0000000000000000000000000000000000,
0000000000000000000000000000000000,
0000000000000000000000000000000000,
0000000000000000000000000000000000,
0000000000000000000000000000000000,
0000000000000000000000000000000000,
0000000000000000000000000000000000,
0000000000000000000000000000000000,
0000000000000000000000000000000000,
0000000000000000000000000000000000,
0000000000000000000000000000000000,
0000000000000000000000000000000000,
0000000000000000000000000000000000,
0000000000000000000000000000000000,
0000000000000000000000000000000000,
0000000000000000000000000000000000,
0000000000000000000000000000000000,
0000000000000000000000000000000000,
0000000000000000000000000000000000,
0000000000000000000000000000000000
);

constant EG_EG_COSH_DETA_LUT_SFIXED : calo_calo_cosh_deta_lut_array := CALO_CALO_COSH_DETA_LUT_SFIXED;
constant EG_TAU_COSH_DETA_LUT_SFIXED : calo_calo_cosh_deta_lut_array := CALO_CALO_COSH_DETA_LUT_SFIXED;
constant EG_JET_COSH_DETA_LUT_SFIXED : calo_calo_cosh_deta_lut_array := CALO_CALO_COSH_DETA_LUT_SFIXED;
constant JET_EG_COSH_DETA_LUT_SFIXED : calo_calo_cosh_deta_lut_array := CALO_CALO_COSH_DETA_LUT_SFIXED;
constant JET_JET_COSH_DETA_LUT_SFIXED : calo_calo_cosh_deta_lut_array := CALO_CALO_COSH_DETA_LUT_SFIXED;
constant JET_TAU_COSH_DETA_LUT_SFIXED : calo_calo_cosh_deta_lut_array := CALO_CALO_COSH_DETA_LUT_SFIXED;
constant TAU_EG_COSH_DETA_LUT_SFIXED : calo_calo_cosh_deta_lut_array := CALO_CALO_COSH_DETA_LUT_SFIXED;
constant TAU_JET_COSH_DETA_LUT_SFIXED : calo_calo_cosh_deta_lut_array := CALO_CALO_COSH_DETA_LUT_SFIXED;
constant TAU_TAU_COSH_DETA_LUT_SFIXED : calo_calo_cosh_deta_lut_array := CALO_CALO_COSH_DETA_LUT_SFIXED;

-- calo-calo cos dphi LUTs
type calo_calo_cos_dphi_lut_array is array (0 to 2**MAX_CALO_PHI_BITS-1) of sfixed(2 downto -19);

constant CALO_CALO_COS_DPHI_LUT_SFIXED : calo_calo_cos_dphi_lut_array := (
010000000000000000000,
001111111110111110011,
001111111011111001110,
001111110110110010001,
001111110000101000111,
001111100111011011001,
001111011101001011110,
001111010000111001010,
001111000010100011110,
001110110010001011010,
001110011111101111100,
001110001100010010011,
001101110110110010001,
001101011111001110110,
001101000110101001111,
001100101100000010000,
001100010000011000100,
001011110010101100000,
001011010011111101111,
001010110100001110010,
001010010010011011101,
001001101111100111011,
001001001011110001101,
001000100101111000110,
000111111111111111111,
000111011001000101101,
000110110001001001101,
000110001000001100010,
000101011110001101010,
000100110100001110010,
000100001001001101110,
000011011101001011110,
000010110010001011010,
000010000110001001001,
000001011001000101101,
000000101101000011100,
000000000000000000000,
111111010010111100011,
111110100110111010010,
111101111001110110110,
111101001101110100101,
111100100010110100001,
111011110110110010001,
111011001011110001101,
111010100001110010101,
111001110111110011101,
111001001110110110010,
111000100110111010010,
110111111111111111111,
110111011010000111001,
110110110100001110010,
110110010000011000100,
110101101101100100010,
110101001011110001101,
110100101100000010000,
110100001101010011111,
110011101111100111011,
110011010011111101111,
110010111001010110000,
110010100000110001001,
110010001001001101110,
110001110011101101100,
110001100000010000011,
110001001101110100101,
110000111101011100001,
110000101111000110101,
110000100010110100001,
110000011000100100110,
110000001111010111000,
110000001001001101110,
110000000100000110001,
110000000001000001100,
110000000000000000000,
110000000001000001100,
110000000100000110001,
110000001001001101110,
110000001111010111000,
110000011000100100110,
110000100010110100001,
110000101111000110101,
110000111101011100001,
110001001101110100101,
110001100000010000011,
110001110011101101100,
110010001001001101110,
110010100000110001001,
110010111001010110000,
110011010011111101111,
110011101111100111011,
110100001101010011111,
110100101100000010000,
110101001011110001101,
110101101101100100010,
110110010000011000100,
110110110100001110010,
110111011010000111001,
110111111111111111111,
111000100110111010010,
111001001110110110010,
111001110111110011101,
111010100001110010101,
111011001011110001101,
111011110110110010001,
111100100010110100001,
111101001101110100101,
111101111001110110110,
111110100110111010010,
111111010010111100011,
000000000000000000000,
000000101101000011100,
000001011001000101101,
000010000110001001001,
000010110010001011010,
000011011101001011110,
000100001001001101110,
000100110100001110010,
000101011110001101010,
000110001000001100010,
000110110001001001101,
000111011001000101101,
000111111111111111111,
001000100101111000110,
001001001011110001101,
001001101111100111011,
001010010010011011101,
001010110100001110010,
001011010011111101111,
001011110010101100000,
001100010000011000100,
001100101100000010000,
001101000110101001111,
001101011111001110110,
001101110110110010001,
001110001100010010011,
001110011111101111100,
001110110010001011010,
001111000010100011110,
001111010000111001010,
001111011101001011110,
001111100111011011001,
001111110000101000111,
001111110110110010001,
001111111011111001110,
001111111110111110011,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000
);

constant EG_EG_COS_DPHI_LUT_SFIXED : calo_calo_cos_dphi_lut_array := CALO_CALO_COS_DPHI_LUT_SFIXED;
constant EG_TAU_COS_DPHI_LUT_SFIXED : calo_calo_cos_dphi_lut_array := CALO_CALO_COS_DPHI_LUT_SFIXED;
constant EG_JET_COS_DPHI_LUT_SFIXED : calo_calo_cos_dphi_lut_array := CALO_CALO_COS_DPHI_LUT_SFIXED;
constant JET_EG_COS_DPHI_LUT_SFIXED : calo_calo_cos_dphi_lut_array := CALO_CALO_COS_DPHI_LUT_SFIXED;
constant JET_JET_COS_DPHI_LUT_SFIXED : calo_calo_cos_dphi_lut_array := CALO_CALO_COS_DPHI_LUT_SFIXED;
constant JET_TAU_COS_DPHI_LUT_SFIXED : calo_calo_cos_dphi_lut_array := CALO_CALO_COS_DPHI_LUT_SFIXED;
constant TAU_EG_COS_DPHI_LUT_SFIXED : calo_calo_cos_dphi_lut_array := CALO_CALO_COS_DPHI_LUT_SFIXED;
constant TAU_JET_COS_DPHI_LUT_SFIXED : calo_calo_cos_dphi_lut_array := CALO_CALO_COS_DPHI_LUT_SFIXED;
constant TAU_TAU_COS_DPHI_LUT_SFIXED : calo_calo_cos_dphi_lut_array := CALO_CALO_COS_DPHI_LUT_SFIXED;

-- muon-muon cosh deta LUTs
type muon_muon_cosh_deta_lut_array is array (0 to 2**(MUON_ETA_HIGH-MUON_ETA_LOW+1)-1) of sfixed(8 downto -19);

constant MU_MU_COSH_DETA_LUT_SFIXED : muon_muon_cosh_deta_lut_array := (
000000010000000000000000000,
000000010000000000000110100,
000000010000000000001101000,
000000010000000000100000110,
000000010000000000111010111,
000000010000000001100010010,
000000010000000010001001101,
000000010000000010111110000,
000000010000000011111001000,
000000010000000100111010100,
000000010000000110000010101,
000000010000000111010111110,
000000010000001000101101000,
000000010000001010001111010,
000000010000001011111000001,
000000010000001101100111101,
000000010000001111100100001,
000000010000010001100000101,
000000010000010011101010010,
000000010000010101111010011,
000000010000011000010001001,
000000010000011010110101000,
000000010000011101011111011,
000000010000100000001001110,
000000010000100011000111111,
000000010000100110000101111,
000000010000101001001010100,
000000010000101100011100010,
000000010000101111110100100,
000000010000110011010011010,
000000010000110110111111010,
000000010000111010110001110,
000000010000111110101010110,
000000010001000010101010011,
000000010001000110110000100,
000000010001001011000011110,
000000010001001111011101100,
000000010001010100000100100,
000000010001011000101011011,
000000010001011101011111011,
000000010001100010011010000,
000000010001100111100001101,
000000010001101100101001010,
000000010001110001111110001,
000000010001110111100000000,
000000010001111101001000011,
000000010010000010110111100,
000000010010001000101101000,
000000010010001110101111101,
000000010010010100111000111,
000000010010011011001000101,
000000010010100001100101100,
000000010010101000001001000,
000000010010101110111001100,
000000010010110101101010000,
000000010010111100101110010,
000000010011000011110010011,
000000010011001011001010010,
000000010011010010100010001,
000000010011011010000111001,
000000010011100001110010101,
000000010011101001101011010,
000000010011110001101010011,
000000010011111001110110110,
000000010100000010001001101,
000000010100001010101001100,
000000010100010011010000000,
000000010100011100000011101,
000000010100100100111101110,
000000010100101110000101000,
000000010100110111010010111,
000000010101000000101101111,
000000010101001010001111010,
000000010101010011111101111,
000000010101011101111001101,
000000010101100111111011111,
000000010101110010000100101,
000000010101111100100001001,
000000010110000111000100001,
000000010110010001101101110,
000000010110011100100100011,
000000010110100111101000001,
000000010110110010111001001,
000000010110111110010000100,
000000010111001001110101001,
000000010111010101100000010,
000000010111100001011111000,
000000010111101101100100010,
000000010111111001110110110,
000000011000000110001111110,
000000011000010010111100011,
000000011000011111101111100,
000000011000101100101111111,
000000011000111001110110110,
000000011001000111010001010,
000000011001010100111000111,
000000011001100010100111000,
000000011001110000100010011,
000000011001111110101010110,
000000011010001101000110110,
000000011010011011101001011,
000000011010101010011001001,
000000011010111001001111011,
000000011011001000011001011,
000000011011010111110000011,
000000011011100111010100100,
000000011011110111000101110,
000000011100000111000100001,
000000011100010111001111101,
000000011100100111101110110,
000000011100111000010100011,
000000011101001001001101110,
000000011101011010001101101,
000000011101101011100001010,
000000011101111101000001111,
000000011110001110101111101,
000000011110100000110001001,
000000011110110010111001001,
000000011111000101010100110,
000000011111011000000100000,
000000011111101010111001111,
000000011111111110000011011,
000000100000010001100000101,
000000100000100101000100011,
000000100000111000111011110,
000000100001001101000110110,
000000100001100001011111000,
000000100001110110000100010,
000000100010001010111101001,
000000100010100000001001110,
000000100010110101100011100,
000000100011001011001010010,
000000100011100001001011010,
000000100011110111011001011,
000000100100001101110100101,
000000100100100100100011101,
000000100100111011100110001,
000000100101010010111100011,
000000100101101010011111101,
000000100110000010010110101,
000000100110011010100001011,
000000100110110010111111101,
000000100111001011110001101,
000000100111100100110000101,
000000100111111110001010000,
000000101000010111110000011,
000000101000110001110001000,
000000101001001011111110110,
000000101001100110100000001,
000000101010000001011011110,
000000101010011100101011000,
000000101010111000001101111,
000000101011010011111101111,
000000101011110000001110101,
000000101100001100101100101,
000000101100101001100100110,
000000101101000110110000100,
000000101101100100001111111,
000000101110000010001001101,
000000101110100000010110111,
000000101110111110110111111,
000000101111011101110011000,
000000101111111101001000011,
000000110000011100110001100,
000000110000111100101110010,
000000110001011101001011110,
000000110001111101111100111,
000000110010011111000001101,
000000110011000000100111010,
000000110011100010100000100,
000000110100000100110100000,
000000110100100111011011001,
000000110101001010100011000,
000000110101101110000101000,
000000110110010001111010111,
000000110110110110010001011,
000000110111011010111011100,
000000111000000000000110100,
000000111000100101101011101,
000000111001001011101011000,
000000111001110010000100101,
000000111010011000111111000,
000000111011000000001101000,
000000111011101000000010011,
000000111100010000001011011,
000000111100111000110101001,
000000111101100001111111110,
000000111110001011100100100,
000000111110110101101010000,
000000111111100000001001110,
000001000000001011001010010,
000001000000110110101011100,
000001000001100010100111000,
000001000010001111001001111,
000001000010111100000110111,
000001000011101001101011010,
000001000100010111101001111,
000001000101000110001001001,
000001000101110101001111110,
000001000110100100110000101,
000001000111010100111000111,
000001001000000101100001111,
000001001000110110101011100,
000001001001101000011100101,
000001001010011010110101000,
000001001011001101100111101,
000001001100000001001000000,
000001001100110101000010110,
000001001101101001101011010,
000001001110011110110100101,
000001001111010100101011110,
000001010000001011000011110,
000001010001000010000011000,
000001010001111001100011000,
000001010010110001110001000,
000001010011101010100110010,
000001010100100100001001011,
000001010101011110001101010,
000001010110011000111111000,
000001010111010100011000001,
000001011000010000011111001,
000001011001001101001101011,
000001011010001010101001100,
000001011011001000110011100,
000001011100000111100100111,
000001011101000111000100001,
000001011110000111010001010,
000001011111001000001100010,
000001100000001001101110100,
000001100001001100000101010,
000001100010001111010000011,
000001100011010011000010111,
000001100100010111101001111,
000001100101011100111110101,
000001100110100011000111111,
000001100111101001111110111,
000001101000110001101010011,
000001101001111010001010011,
000001101011000011011000010,
000001101100001101100001000,
000001101101011000010111110,
000001101110100100000010110,
000001101111110000101000111,
000001110000111110000011011,
000001110010001100010010011,
000001110011011011011100010,
000001110100101011011010101,
000001110101111100010100000,
000001110111001110001000011,
000001111000100000110001001,
000001111001110100011011011,
000001111011001000111010001,
000001111100011110010011110,
000001111101110100101111000,
000001111111001100000101010,
000010000000100100010110100,
000010000001111101101001010,
000010000011010111111101100,
000010000100110011001100110,
000010000110001111011101100,
000010000111101100101111111,
000010001001001010111101001,
000010001010101010011001001,
000010001100001010110000001,
000010001101101100001111001,
000010001111001110101111101,
000010010000110010010001110,
000010010010010111000010100,
000010010011111100110100110,
000010010101100011101111001,
000010010111001011111000001,
000010011000110101000010110,
000010011010011111011011111,
000010011100001010111101001,
000010011101110111101101001,
000010011111100101100101001,
000010100001010100101011110,
000010100011000101000001001,
000010100100110110100101000,
000010100110101001011110001,
000010101000011101011111011,
000010101010010010110101110,
000010101100001001100001011,
000010101110000001011011110,
000010101111111010110001110,
000010110001110101010110011,
000010110011110001010000010,
000010110101101110100101111,
000010110111101101010000101,
000010111001101101010111001,
000010111011101110110010111,
000010111101110001101010011,
000010111111110110000100010,
000011000001111011110011010,
000011000100000011000100100,
000011000110001011111000001,
000011001000010110000001000,
000011001010100001110010101,
000011001100101111000110101,
000011001110111101111100111,
000011010001001110010101100,
000011010011100000010110111,
000011010101110011111010101,
000011011000001001000111010,
000011011010011111111100101,
000011011100111000100001100,
000011011111010010101000110,
000011100001101110011111010,
000011100100001100000101010,
000011100110101011011010101,
000011101001001100011000111,
000011101011101111001101001,
000011101110010011110000110,
000011110000111010001010011,
000011110011100010011010000,
000011110110001100011111100,
000011111000111000011011000,
000011111011100110001100011,
000011111110010101111010011,
000100000001000111100100111,
000100000011111011001011111,
000100000110110000101111100,
000100001001101000001111100,
000100001100100001110010101,
000100001111011101011000111,
000100010010011011000010001,
000100010101011010101110011,
000100011000011100100100011,
000100011011100000011101011,
000100011110100110100110101,
000100100001101110110010111,
000100100100111001001111011,
000100101000000101111100000,
000100101011010100110010011,
000100101110100101111111011,
000100110001111001011100100,
000100110101001111010000011,
000100111000100111010100100,
000100111100000001110101111,
000100111111011110101110000,
000101000010111101111100111,
000101000110011111101111100,
000101001010000011111111100,
000101001101101010101100110,
000101010001010011110111011,
000101010100111111101100010,
000101011000101110000101000,
000101011100011111000001101,
000101100000010010101000110,
000101100100001000111010001,
000101101000000001110101111,
000101101011111101100010101,
000101101111111100000000011,
000101110011111101001111000,
000101111000000001010101001,
000101111100001000001100010,
000110000000010010000001011,
000110000100011110101110000,
000110001000101110010010001,
000110001101000000111010111,
000110010001010110100001110,
000110010101101111001101001,
000110011010001010110110101,
000110011110101001101011010,
000110100011001011101011000,
000110100111110000110110000,
000110101100011001000101101,
000110110001000100101101011,
000110110101110011100111000,
000110111010100101110010010,
000110111111011011001111010,
000111000100010100001011000,
000111001001010000011111001,
000111001110010000010010000,
000111010011010011100011101,
000111011000011010011010110,
000111011101100100110111010,
000111100010110010111001001,
000111101000000100100000010,
000111101101011001111010000,
000111110010110010111111101,
000111111000001111110111110,
000111111101110000100010011,
001000000011010101000110000,
001000001000111101100010101,
001000001110101001111110111,
001000010100011010010100010,
001000011010001110101111101,
001000100000000111010001010,
001000100110000011111001000,
001000101100000100100110111,
001000110010001001101000000,
001000111000010010110101110,
001000111110100000010110111,
001001000100110010010001110,
001001001011001000011111111,
001001010001100011001110011,
001001011000000010011101010,
001001011110100110001100011,
001001100101001110100010100,
001001101011111011100110001,
001001110010101101010000101,
001001111001100011101111001,
001010000000011110111011001,
001010000111011111000001101,
001010001110100011111100010,
001010010101101101111000000,
001010011100111100110100110,
001010100100010000110010110,
001010101011101001111000011,
001010110011001000001100010,
001010111010101011101110011,
001011000010010100100101010,
001011001010000010101010011,
001011010001110110010001011,
001011011001101111010011110,
001011100001101101111000000,
001011101001110001111110001,
001011110001111011101100101,
001011111010001011010000111,
001100000010100000011101011,
001100001010111011100110001,
001100010011011100100100011,
001100011100000011011110110,
001100100100110000011011110,
001100101101100011100010000,
001100110110011100101011000,
001100111111011100001010001,
001101001000100001111001001,
001101010001101101111110100,
001101011011000000100000110,
001101100100011001011111110,
001101101101111001001000111,
001101110111011111011011111,
001110000001001100011000111,
001110001011000000000110100,
001110010100111010110001110,
001110011110111100010100000,
001110101001000100111010100,
001110110011010100100101010,
001110111101101011011010101,
001111001000001001011010111,
001111010010101110111001100,
001111011101011011110000000,
001111101000001111111110010,
001111110011001011111000001,
001111111110001111011101100,
010000001001011010101110011,
010000010100101101110001011,
010000100000001000110011100,
010000101011101011110100111,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000,
000000000000000000000000000
);

-- muon-muon cos dphi LUTs
type muon_muon_cos_dphi_lut_array is array (0 to 2**(MUON_PHI_HIGH-MUON_PHI_LOW+1)-1) of sfixed(2 downto -19);

constant MU_MU_COS_DPHI_LUT_SFIXED : muon_muon_cos_dphi_lut_array := (
010000000000000000000,
001111111111111001011,
001111111111110010111,
001111111111011111001,
001111111110111110011,
001111111110011101101,
001111111101110110010,
001111111101000001111,
001111111100000110111,
001111111011000101011,
001111111001111101010,
001111111000101000001,
001111110111001100011,
001111110101110000101,
001111110100000111110,
001111110010010001110,
001111110000011011110,
001111101110011111010,
001111101100010101101,
001111101010000101100,
001111100111101110110,
001111100101010001100,
001111100010100111000,
001111011111111100101,
001111011101000101001,
001111011010000111001,
001111010111000010100,
001111010011110111011,
001111010000100101101,
001111001101001101011,
001111001001101000000,
001111000110000010101,
001111000010010000001,
001110111110010111001,
001110111010010111100,
001110110110010001011,
001110110010000100101,
001110101101110001011,
001110101001010001000,
001110100100110000101,
001110100000000011010,
001110011011001111010,
001110010110011011001,
001110010001011010000,
001110001100010010011,
001110000111000100001,
001110000001101111011,
001101111100010100000,
001101110110110010001,
001101110001001001101,
001101101011011010101,
001101100101100101001,
001101011111101001000,
001101011001100110011,
001101010011011101001,
001101001101001101011,
001101000110110111000,
001101000000010011101,
001100111001110000001,
001100110011000110001,
001100101100011100010,
001100100101100101001,
001100011110100111100,
001100010111100011010,
001100010000011000100,
001100001001001101110,
001100000001110101111,
001011111010011110000,
001011110010111111101,
001011101011011010101,
001011100011101111001,
001011011011111101001,
001011010100000100100,
001011001100001011111,
001011000100000110001,
001010111100000000011,
001010110011110100000,
001010101011100001010,
001010100011000111111,
001010011010101110011,
001010010010001110100,
001010001001101000000,
001010000000111010111,
001001111000001101111,
001001101111011010010,
001001100110100000001,
001001011101011111011,
001001010100011110101,
001001001011010111011,
001001000010001001101,
001000111000111011110,
001000101111100111011,
001000100110001100011,
001000011100110001100,
001000010011010000000,
001000001001101000000,
000111111111111111111,
000111110110010001011,
000111101100100010110,
000111100010101101101,
000111011000110001111,
000111001110110110010,
000111000100111010100,
000110111010111000010,
000110110000101111100,
000110100110100110101,
000110011100010111010,
000110010010000111111,
000110000111111000101,
000101111101100010101,
000101110011000110001,
000101101000110000010,
000101011110001101010,
000101010011101010010,
000101001001000111010,
000100111110100100001,
000100110011111010101,
000100101001010001000,
000100011110100000111,
000100010011110000110,
000100001001000000101,
000011111110010000100,
000011110011011001111,
000011101000100011001,
000011011101100101111,
000011010010101111010,
000011000111110010000,
000010111100110100110,
000010110001110001000,
000010100110110011110,
000010011011110000000,
000010010000101100001,
000010000101101000011,
000001111010100100101,
000001101111100000110,
000001100100010110100,
000001011001010010101,
000001001110001000011,
000001000010111110000,
000000110111110011101,
000000101100101001010,
000000100001011111000,
000000010110010100101,
000000001011001010010,
000000000000000000000,
100000001011001010010,
100000010110010100101,
100000100001011111000,
100000101100101001010,
100000110111110011101,
100001000010111110000,
100001001110001000011,
100001011001010010101,
100001100100010110100,
100001101111100000110,
100001111010100100101,
100010000101101000011,
100010010000101100001,
100010011011110000000,
100010100110110011110,
100010110001110001000,
100010111100110100110,
100011000111110010000,
100011010010101111010,
100011011101100101111,
100011101000100011001,
100011110011011001111,
100011111110010000100,
100100001001000000101,
100100010011110000110,
100100011110100000111,
100100101001010001000,
100100110011111010101,
100100111110100100001,
100101001001000111010,
100101010011101010010,
100101011110001101010,
100101101000110000010,
100101110011000110001,
100101111101100010101,
100110000111111000101,
100110010010000111111,
100110011100010111010,
100110100110100110101,
100110110000101111100,
100110111010111000010,
100111000100111010100,
100111001110110110010,
100111011000110001111,
100111100010101101101,
100111101100100010110,
100111110110010001011,
100111111111111111111,
101000001001101000000,
101000010011010000000,
101000011100110001100,
101000100110001100011,
101000101111100111011,
101000111000111011110,
101001000010001001101,
101001001011010111011,
101001010100011110101,
101001011101011111011,
101001100110100000001,
101001101111011010010,
101001111000001101111,
101010000000111010111,
101010001001101000000,
101010010010001110100,
101010011010101110011,
101010100011000111111,
101010101011100001010,
101010110011110100000,
101010111100000000011,
101011000100000110001,
101011001100001011111,
101011010100000100100,
101011011011111101001,
101011100011101111001,
101011101011011010101,
101011110010111111101,
101011111010011110000,
101100000001110101111,
101100001001001101110,
101100010000011000100,
101100010111100011010,
101100011110100111100,
101100100101100101001,
101100101100011100010,
101100110011000110001,
101100111001110000001,
101101000000010011101,
101101000110110111000,
101101001101001101011,
101101010011011101001,
101101011001100110011,
101101011111101001000,
101101100101100101001,
101101101011011010101,
101101110001001001101,
101101110110110010001,
101101111100010100000,
101110000001101111011,
101110000111000100001,
101110001100010010011,
101110010001011010000,
101110010110011011001,
101110011011001111010,
101110100000000011010,
101110100100110000101,
101110101001010001000,
101110101101110001011,
101110110010000100101,
101110110110010001011,
101110111010010111100,
101110111110010111001,
101111000010010000001,
101111000110000010101,
101111001001101000000,
101111001101001101011,
101111010000100101101,
101111010011110111011,
101111010111000010100,
101111011010000111001,
101111011101000101001,
101111011111111100101,
101111100010100111000,
101111100101010001100,
101111100111101110110,
101111101010000101100,
101111101100010101101,
101111101110011111010,
101111110000011011110,
101111110010010001110,
101111110100000111110,
101111110101110000101,
101111110111001100011,
101111111000101000001,
101111111001111101010,
101111111011000101011,
101111111100000110111,
101111111101000001111,
101111111101110110010,
101111111110011101101,
101111111110111110011,
101111111111011111001,
101111111111110010111,
101111111111111001011,
110000000000000000000,
101111111111111001011,
101111111111110010111,
101111111111011111001,
101111111110111110011,
101111111110011101101,
101111111101110110010,
101111111101000001111,
101111111100000110111,
101111111011000101011,
101111111001111101010,
101111111000101000001,
101111110111001100011,
101111110101110000101,
101111110100000111110,
101111110010010001110,
101111110000011011110,
101111101110011111010,
101111101100010101101,
101111101010000101100,
101111100111101110110,
101111100101010001100,
101111100010100111000,
101111011111111100101,
101111011101000101001,
101111011010000111001,
101111010111000010100,
101111010011110111011,
101111010000100101101,
101111001101001101011,
101111001001101000000,
101111000110000010101,
101111000010010000001,
101110111110010111001,
101110111010010111100,
101110110110010001011,
101110110010000100101,
101110101101110001011,
101110101001010001000,
101110100100110000101,
101110100000000011010,
101110011011001111010,
101110010110011011001,
101110010001011010000,
101110001100010010011,
101110000111000100001,
101110000001101111011,
101101111100010100000,
101101110110110010001,
101101110001001001101,
101101101011011010101,
101101100101100101001,
101101011111101001000,
101101011001100110011,
101101010011011101001,
101101001101001101011,
101101000110110111000,
101101000000010011101,
101100111001110000001,
101100110011000110001,
101100101100011100010,
101100100101100101001,
101100011110100111100,
101100010111100011010,
101100010000011000100,
101100001001001101110,
101100000001110101111,
101011111010011110000,
101011110010111111101,
101011101011011010101,
101011100011101111001,
101011011011111101001,
101011010100000100100,
101011001100001011111,
101011000100000110001,
101010111100000000011,
101010110011110100000,
101010101011100001010,
101010100011000111111,
101010011010101110011,
101010010010001110100,
101010001001101000000,
101010000000111010111,
101001111000001101111,
101001101111011010010,
101001100110100000001,
101001011101011111011,
101001010100011110101,
101001001011010111011,
101001000010001001101,
101000111000111011110,
101000101111100111011,
101000100110001100011,
101000011100110001100,
101000010011010000000,
101000001001101000000,
100111111111111111111,
100111110110010001011,
100111101100100010110,
100111100010101101101,
100111011000110001111,
100111001110110110010,
100111000100111010100,
100110111010111000010,
100110110000101111100,
100110100110100110101,
100110011100010111010,
100110010010000111111,
100110000111111000101,
100101111101100010101,
100101110011000110001,
100101101000110000010,
100101011110001101010,
100101010011101010010,
100101001001000111010,
100100111110100100001,
100100110011111010101,
100100101001010001000,
100100011110100000111,
100100010011110000110,
100100001001000000101,
100011111110010000100,
100011110011011001111,
100011101000100011001,
100011011101100101111,
100011010010101111010,
100011000111110010000,
100010111100110100110,
100010110001110001000,
100010100110110011110,
100010011011110000000,
100010010000101100001,
100010000101101000011,
100001111010100100101,
100001101111100000110,
100001100100010110100,
100001011001010010101,
100001001110001000011,
100001000010111110000,
100000110111110011101,
100000101100101001010,
100000100001011111000,
100000010110010100101,
100000001011001010010,
000000000000000000000,
000000001011001010010,
000000010110010100101,
000000100001011111000,
000000101100101001010,
000000110111110011101,
000001000010111110000,
000001001110001000011,
000001011001010010101,
000001100100010110100,
000001101111100000110,
000001111010100100101,
000010000101101000011,
000010010000101100001,
000010011011110000000,
000010100110110011110,
000010110001110001000,
000010111100110100110,
000011000111110010000,
000011010010101111010,
000011011101100101111,
000011101000100011001,
000011110011011001111,
000011111110010000100,
000100001001000000101,
000100010011110000110,
000100011110100000111,
000100101001010001000,
000100110011111010101,
000100111110100100001,
000101001001000111010,
000101010011101010010,
000101011110001101010,
000101101000110000010,
000101110011000110001,
000101111101100010101,
000110000111111000101,
000110010010000111111,
000110011100010111010,
000110100110100110101,
000110110000101111100,
000110111010111000010,
000111000100111010100,
000111001110110110010,
000111011000110001111,
000111100010101101101,
000111101100100010110,
000111110110010001011,
000111111111111111111,
001000001001101000000,
001000010011010000000,
001000011100110001100,
001000100110001100011,
001000101111100111011,
001000111000111011110,
001001000010001001101,
001001001011010111011,
001001010100011110101,
001001011101011111011,
001001100110100000001,
001001101111011010010,
001001111000001101111,
001010000000111010111,
001010001001101000000,
001010010010001110100,
001010011010101110011,
001010100011000111111,
001010101011100001010,
001010110011110100000,
001010111100000000011,
001011000100000110001,
001011001100001011111,
001011010100000100100,
001011011011111101001,
001011100011101111001,
001011101011011010101,
001011110010111111101,
001011111010011110000,
001100000001110101111,
001100001001001101110,
001100010000011000100,
001100010111100011010,
001100011110100111100,
001100100101100101001,
001100101100011100010,
001100110011000110001,
001100111001110000001,
001101000000010011101,
001101000110110111000,
001101001101001101011,
001101010011011101001,
001101011001100110011,
001101011111101001000,
001101100101100101001,
001101101011011010101,
001101110001001001101,
001101110110110010001,
001101111100010100000,
001110000001101111011,
001110000111000100001,
001110001100010010011,
001110010001011010000,
001110010110011011001,
001110011011001111010,
001110100000000011010,
001110100100110000101,
001110101001010001000,
001110101101110001011,
001110110010000100101,
001110110110010001011,
001110111010010111100,
001110111110010111001,
001111000010010000001,
001111000110000010101,
001111001001101000000,
001111001101001101011,
001111010000100101101,
001111010011110111011,
001111010111000010100,
001111011010000111001,
001111011101000101001,
001111011111111100101,
001111100010100111000,
001111100101010001100,
001111100111101110110,
001111101010000101100,
001111101100010101101,
001111101110011111010,
001111110000011011110,
001111110010010001110,
001111110100000111110,
001111110101110000101,
001111110111001100011,
001111111000101000001,
001111111001111101010,
001111111011000101011,
001111111100000110111,
001111111101000001111,
001111111101110110010,
001111111110011101101,
001111111110111110011,
001111111111011111001,
001111111111110010111,
001111111111111001011,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000,
000000000000000000000
);

end package;
