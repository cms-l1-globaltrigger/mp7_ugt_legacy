-- Description:
-- Package for LUTS with sfixed format values.

-- Version history:
-- HB 2020-03-14: first design

library ieee;
use ieee.std_logic_1164.all;
-- use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
-- use ieee.numeric_std.all;
use ieee.fixed_pkg.all;

-- use work.lhc_data_pkg.all;
-- use work.math_pkg.all;
use work.gtl_pkg.all;

package sfixed_luts_pkg is

